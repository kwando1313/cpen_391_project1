��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�6�!�~�\@NQzB5�1�kR8�W��7�����e6� �����ْ����5�}܇��M� f�/�_�p���Y۪�^�ow��PS�*'��,e�/�W^j��������ք��ݜQRiZ�-
�}u�d�|"4�����fTD~e{�I��ks�W�oKG��]��6Du������V���r@�Wcle5�t��"��a�ǎ����"b:ٯ��O�A���k���֩y
�^P��}cC5	,R�W)��ɑ"�C��Wh9U�sɕ�B{�T��'���Ч�k/Ƭ��7�kֳ�q��	�c8Y�&s�mCM���lZ�~>�f7@��(�a�JL/��������Ly���C�2g�& ;���ս�\w���Hu���4J4Y���!P*Z_|޼��1xA�/���m�������/&���Cʿ(
��,@�d܈�K����~?8�d���s�s��c�8܂��l���SX��G2�`�<Tt5iP&JP�2�8|�1*�)юa��А�t������p���������7?}�s�{��־���l����M}�)� _
�o��&pPW>���X+R�T��<�V������4�\-N�����U�g H3$#6
�q�֕�,Wz}��E��ۅ��Zdc��(���f�6 "4����a�O̀�R�mrM��?��Cgh��7L�����43K�ե��Ƈ���3ylc���}�Ū�`O��b��R�|t�����.���!�F#�0�}.*:"���|�����Z:E�\�d�I�\Q0����v�֯w�j����Ć,{�+b�Q~�X0�h�(D���p;蜁�!p+~MP�O��X#-t��f}Ɏo��`R>V>�����^��]W�X$�7ˀ����KҚڥ�}��7�����*�דyRQ��#[�H"Q+���A�ÿD{�@�
��LH=֜B_�,g�B@P�S*�[f�y�1�+b������N��l�e(<B��R����(�yu�)��?����O]��EW���(jʄ��t��G���K��EӮf��_�E��vQO�e�ƻ��mՀe��L$�$�=���dr�:�Ru��lJ�]��Ʃ+Q�T��ڙr.*��]C�^Eewt\^.�}zd:=s�tuy�1}��j6<��m�U{�G�|ګ������˺2f��z	��w_8%��(�ŗ^��^�Q�rN3����A�~���h���z��9��f�sp�������B�8���ڷD�'���Л�5,쀟�M�
fZy` "��C�k�>���M4i��S�@�s���%��w�?�L�t��Ġ�0Wb���B�G�#�X�ٵ-�M;xd�Ē�	!6A��K���1����7]:j��BP`�FF",ǘ��_��{�0ֱ/�H^6�,�2�'�ER����9*!��F�uh��m�%�A�LY�X����V���O�
Y�g@����ưl�/�Je%�y1B��~p1�!�b��L�h���b�QF�.���B�/$��G`Or0�%��婺�v֠#��X�gW�Kru��V��-��Q�&�i]�-O�w�8梀l�$Շ|f�F�� o���!���t�Yk��U/D�8��v��L&�w$��(@a:��+��������!&��r�h{����P��cV*�{o��[t�m��Y�0�r0͠�#��g��j�;��[OWd6v$$�1�]��PJ$�0YY����p�['dȒH�Z N�[I�� Kw��m�
͌.u�6�:g���(�����"\X�9I�y��B��'��$�Ā��"%G�Zm�'�A�kYsBH� zrz�����]�+�:ូn9z��G	���u{�.v&=����Qia-��)Y�u�	�LZ|ct�� S���#�|�k��H!�鳛Ǉ;йs�}z`��1G)�);�	�א��T��kl�ϣ,����j�a���6l/}���M��+I5 �����  �=�f[R#Z/�{s��~n�y��eT(��t���Q2���O���K���`2P�w��@Am��wD��Vd�@��_!�B��F�$}i�O<�& �B>/��㴹	���1eu��]f@�CI��W�"���ofc7f��@B�tU���e�.��:�������o�ϓ�^���~&�k�DZ�l���M�8��<���t��[3�i�
�{8<�\^at��V����}�A��,d-�h�n���4�{n�U�q	��:�4F����(!�����vJf���e�R91a��#�d\&�z�1��#!�f��!�g2d�Hwc�ц]���S�ުz3H>��C�F���S�����a�œcBԻĤni_/9yA��`�9��;W�E���9���v��=ꭖZ'�uo<�kd�Ɓ+7�u
��S����w^��9ݢd6p�L�m��l�U��3֐/�h�i��#�����\�C�����BZƬgAŇ;�F&���Q~*Y�JQ�R`�&'���wѾ� IL�rQS��|?՘�s3P���}+<m�rq�೩���	 Q�RXX�F���������&���_�/���h�����}�t����ݣ���]u��J��i����j!_`U�<as���'��+sҵ��5"��p�	��:�ؾX>1U�u�86u6Q���p33�������̋u ^P*�9�JN�ӝ�<���>8��?;��R�n7��Q_HJ��P1t��jI��*��]�H�_b�<v������(ͧc�U��ꝶ�|K=�����6���T�0:`�dd����Hn� �W	P�7w�$O��;T�;��|}́jSܼ�n�!2���d�w8޷���&^K�=.(��]�~Sa�	��>�JI�k6c�yt^�J�����B{rF\j��x(,�4ǒ����Ҕ��#ހl�y�k}~+yX2�h.�7��2˸͙we���V4r�u�;�R=��$�q��,�j�ܓcU�kyv�Y=�*�^]bYD4��͓�^m\�F�s�+���I2�'��+��Yq��#�2���S�Jg��Aj�Py
"6��>Ƒ�����f�"�!5dŷ�*e�|�):-�z����ǀN�e�̹�<�vKe_Mޝ3:$}&�1�R��I4ϒ�N����oe,�%�6}�m���j�7mP(� �����Ć��=�i��uq=�5
���{�|f�k:������N;��"�r�Q;߶��]a~�e�4�7MY>�7�!�|�GO��0�-�Z�(U!��ِY��h�
b�Q�%9NB�� R��2��J�@a�^�w8�}�QUF!B��C�J(�v������{+m,�M�:�d���ܽal��۸�|�^����� L|M9D�Y-��op\�����4����75 ���kiO&�/���ʭ�7�=��,zآ�We�.p�o��kJ��R��T�^�����^D,��iS�|UV�Djm�e���ͽ��0���|��}M���J��	oM�c�s��=>�a�f$@��7���RgJ�y�T�	�P��9�{Mg�r��r^(�
��lq��e;	c镢�YΈ���-�
�ݥ���<,]���6Xm��"y�+ĩz}�C��Uj�;�*4<����o��"���UH��^(\�u�i�Y|Z�so\��*�8�����j�7�1/�`��x6#+C��Ъ��K�����;�n��	���s/xo���37�q��Hs��6|�_�ȉ�#\��?��a�N�֍��/*M�
��R��Ák���"�M�B�.���m#�o��4�(u�Q2q��Yf�D`@��Kimb�Ц}&꓇}���#ava�?q��(6�([�}���x���÷H���Y��x'd�e�KWǱUj��8]4' 얹>+��>�	V��q�X�`��g+hcg���}v9�|��W���g�j���Uc����d��T"	F�H�d7�=X����.ͥY��^�;7��n���[ǩFU���/5 v�d�=IX܉s^�r@~�'m��QW�$�7_Bҫ'��$�7	(��!C�8\�Ï-f.K�d.DE}W0hB��7�X�p�v��C����R�q�d�@�a8������P�Q޻�H�UT5v��jm��\�\hל�I��a�%	���a3��d�`h8\�V�
�(�����Z�(��
����+��wc�Z�'���		U��N��n&wK:��D��
�lO0X���5��(L���r�I���bGY��U��N�6@��O|��]z���&�m�!��̩�S�*�����$"w�@C�����h5�^T�?�$hh��<����;@�N���ĥc�����8ϑ��j�<
A~��,�u.�� �-�]�.��,)��g\��Y<� �<�b��=
�nf�|�n`����ضm��a;�`�:z��D�ѓ��a2)�ұ�����۱�;��_n{��X=�:%��q���լ�}j�x@r�--E����c"<��}	��M���3ZwUIR����wg��AHV�o��I�u�u�|7@X�A@����D:O>j����c��L�����zЍI3�����<8����/��~x(]��j$���j�&)u/}��X���j�.����ab얶���TN�;����dxT��n���#�,p{�{���Q�?LsU�� � �B�y���9 �����E�*����N���q8�0]Bݖ��]	I5Kh6+|�9Y�[,�Q�u;s��g�Q��z�W��j������gS���{���1�K5�ajBH�&�k�Ӕ,�˝���ԨY!n�Ta�^�N�E֡��V|�{�$$�f�+wu���E�"���>@ɿ�sh�SLH]<���1롮�E"�ht�Δ�l�����4��da�k��ߴ��v�q��gQn�-O�Ɓ;��%�\�g�3(9�Yx� �����I1�	h�W=�|¤�j�U��D��L�G���bـ�n ��"��9�o�O/��LP٪��"n��ޭ��ؾ@0ԋ	A6;�����lZ��͒8T����Ղ�$�Ag��R��x=4��+�>g�=��u칓Ԡ�ݜ' �}z+EW�ܝɊ�Lv��ލ���' ��y��<�_���S���vz�����+W�H#���Y�[m�N#bpj��2��<D�'�T1z�i�h�j�1�w�\sW���"�Ƌ�hɖ�܅ߢf��tm�v�n�L�j�/�k,B��֑QȤ�0>ԝ>A��fۀ���,�e��h�T/b�����Π����-��@��D����3$����BŒnx��)�����ߡ�F*)�4����X^̱"ds���Ѳ��ј�F&ޞ��CW� �2�[��̅:D֪��
�ߠe�OT|H�t�5���']�ٖX!s�A�b��p��
��.dZ�H��do"�m평����|Z)�E�1D�O�[��ZmE@ʎJ���̽����&c;ܧ��6 t�|�����E�O�ELu��JɈ�S�b�(��� gA������@�U��P$�)�4�f׏��rݥ�&&�j�~�X���_w6�J�iď2k5K�d笠���t���V�/��A�d���ѫ[[�n9P���^Ք$`�B}�If���@����p�Ǒ��%�Ħ�+�qҷ�.��:љcpR��uab:~��@r¨��7gS�a�l�������!&�P��55�a��]����s��+jʽ�H��v�3�����hD��0�:I	�g�����DNZ$f:��T��`��\��c�Z����?/�$�c��Xf��O���e�ԮT8\�-��k�p5|�\\V��??-��o
4Q��M&G�䵈�'=|	T��HDN!w�����<i��Wx$mV�_���n��]z��i�J��TV�ɮh�y���.�/z�-ng��h�0�y��&1,UVF7�1߀0�F51��w��R�70,���DҠ
��6LS\v�X��Ab]�~!��1W��Z�6d{)u�~��_!ދ��]�Vt���76,��?��k7�2@R�*���%rW����KX�4�{��b�lĿ:����g�ԟl"�}0x넢��F�))�*��<�4!6u���L��7mQ�T�18��(B���~?S�o�&��-d�����`
 �H�ʦ�q�l!��qtV����Zn�����ǡVzb�:�ҫ<�n|�g��Kٳ��@�)�|9���v���dݽ{������I>��@�4N�sǯ!2���_}]� ^���[qr�����,��.���46�ʽ��
�XBǍ�Y-��-��F=�^�����w�hH��>���1�Ұ��j��a+T���&ߜ������7����
=d���������=5�@b*��f��]T��q������������j�5$�S�IC���g-�xn��)�ݺ�����#u��%)'�Ϧ�Hu�������!7xHc�=����}-{����yo��_�J '���V���`:
c�-��e�������BR�=XB�<)����K�:����sufElS������'&�Ш�f�Y���m���P민�]�7�Z}Aɹ�w�.���'�ewz.H�YC�5�,�����Q�uҦoք�D���յ�����O"�� �aoVv��|ǘӁ��(��t���u���?wGpn�6w1�pTI`q7��#F؈�=��W��%N��Z�:b]&�9��C#Ш]���L�˗����1�����"�l���vi�ӳ_��;l��o.��x�l���_�>�|����d���`PlG�zGA7���+��~h���$��������̾�q��j�Wۢ���O䁀(���+Vƹ�v���- X�N��9��>�.x4����E����et>���*1ѝb�dT������w��}T�p����.�(�R��S�<f�@h�<;K��o��8�,�k
+��J@�TEn��K�,ܡ��C�]MR�JpHji�ְ��jb!K{�V�U�Vx��Ԅ@y>D@����$1鋤P��Z�������8Bg���x�\t��"����5ޅ�6��#0MC�Q����z�P����C�9�=����L-H�S{���gd�m�8�X3��f�.@�\�K�|�W�$�o9j���ϸѸ\�ooGT2G,^
��}�|�{���4KZ���a�6X�#H�@:�g��.�Lz[�{�1���%�ޫ �j@�s������mI::��Fr$���ty�����w���k|�3��x��Wp��;�K(���'��gqtϷ��L䭠	$��g��Wk�{�+LS#ڑ��AV�_I��J�4�@���L�����sG�!0���Q�fU����oQ|=Ъ���1��=#N��B���ʜ�%R�UXz8��%�
���W;.�ʨ�Hb�$7x�g}���AL��S�يͽ���)ͻ��6����*r��/���y�sɳe�wv���t��y���>ù�Ÿ���E�D�;�O �n�a�ZČ	[�Ο݈cz�q��ᅴm��"�@����[~�E}�R@���l�O���u�uH��VY���;k������ڲC"ᤊvP�-0��ZjvU;��
�u�w�d�Zުo �^�t&���st�5��t�"0�#�s#t�h����z��b�(���P١���d���NwbV�!;���f��D�/alXm�d�HV��]��+5���� �B4�{Mh��hf54��)��Kf��0Zu�<���A�2{Y��#T`%�U#���/��P�--��Q�O��
W���,!�%[���Ty�հWNQצ�LC2A�G�-UA�-B�2���}�� ��h�C�R��)<h�<�]�S�F��;|��5���P/	���]��ߔg=�����7��@�6�|x���i�����k.�\c�f#�,�X�(ԛR݉3�5Fg^���������jA|*�M֏���'=��hم�ղ��^7;��g�e�hI� 2L��7���kQ�^۬#�ї��M_�IGr����ŊF(Pջ�������L9��4F-)��{�.k�8�Ř){�SJ�\�?�S���b�L�O�ᢦ�A0���� �(��ͧ��e�~%�����pV�[���J��8h�~�^�k���gC���N�����>J!�v�����ݡ�H����BM���WZ�g�\���"�z�0U�G.��j[� �rp%gH�FN���9�,o¿�1�y�j��q�Ky����O��@:��������+;8kT.���g����d�}��R"��n+�5�����|��ػ$䪪�#�xT����m����Z7���s	���� zX��Lc_����<�^]���`�K��{�<z�y��N
վ��:e'U}fm��]��`&�!�%֐�V���R`�'c'Ӏ��}���e3���c�7�bcw�N�C3)����s�:�jO�,��A��;��ٞx8;�}��CFUy�F�(v��h�Y�v����`�}�v��CkUh�#gү��|O����n;'���n��8���ʄ���ګ�B/�妨(��F����r���Gm���a]��2���"�E�����4��&�s>��F��T=�G�x�5C����+s��-��i��N�0
H��fo�9k����ʠ-@�խ��(S���'/�C��%��jn

���@���Q��8D ����C��J�k�;������K��p~�p"�x�~�c��²�����j��C�UŹV/�(|u��O\�������yPf���L��O���-M��>>�L�<IZ>��C�\��a��8�"��4W����b�e�'�h�� ��p�<>�7+$P��wx2[L|��~�
q���V�|���$� �5�1�Q�?��J�$�T�
�'��i3>6|�RA��{c��G���B���1o1�*�
B����Us��� ���@��:�K�6��K�m9!�P�Eq�
gtǲ~49r���@r�
��,�A�����������7�rg4r�'^ڽ��D��J�����փ�����7��&��W�\�ؒ�jE�Q�SNۧ%�8]�� scb��Z�����c2���6��~�f���̺�w-\L����7��\��њ�p�XCȁ����fZ0���7 ���7Q�R����U�mI������
_�c,�xQ�$Ûp���H�E�=�*Y�4��=P9�@��G�	�����ڟLW!%8J�F5����b��c��t���\���]�T��	YIl��%�,�;΃$��.-
M�1u�}$��?`���*�>hdj,��uM �T���|��?Sv!��E�Ƣb�Fu�)=���Vۯ�L�Y���*�MªUu��g�j�uk'%�{�-b�e�~�vނ�7S:T���w��vE_�) ���Bp]��T��\�^�L��m��S���o#������.����3v�s@�T���#P̹�W��U�%�簹zG��,":Կ�l�����D>��v��F�5�\q�X�x����������Pc]�/� ����'4Y*��f�0m�qR���u�a������y$��e�>^ˊ�
@㝖aU��FeG����RB�a9�&��{��C]��63P�x��kM�5��=a��מ(uK@��j3�!����5b���g�#N~��o�1���2����×��B#��^+m��2jЬ	��(�$4��[N�I����K��5�����e����˱��"�62ͬF9���Kk���1ߞ�'D� Y��i��E�k|��t��S�^��t>zz��!}�����p�����P��Do���f^R�u���ҝv;�},<>}���_�IiC
�ħ�TF��Po��'��2�x�0�>�(������Oሠ��"\��6ܹ�u%��$taЄ�!١�V��/:I��z�e`� D��`�5~�P�4oŒ�����pm�K��K8T�ƹ܎x�ӫ��!��mD��v����_�b��A��]S�/��O�w/�%��F��	�x���\�+b5>8�9��#�y�q�_�=ٹ�xr���vmɂ���!���b��1>gM������ ��R�d֌	����t�h;ر�i�-�y��8=w�U�<�s���&#�Ok����̔�:l�ޣ�z� (��+�'y�?�����O��G�mV���1H�p�}����{\w�	���[ BBٛ�f�2*T�#���W5���_V�a���� �;S��j�����)��Y vQ"�OJ�!^őBl W��E�LU�|5(�|�Y1���O��/���5�+ZI~wz�*��a'��|b,��
m�����x�#AVu��%�Õ{���E7�U��q%&dKZ�ƙ:��B��0�o3=Xǐ�D��p㵈�%�+�̜��W����ۙ����y�����}�P{��oE�txq���Hox���ü����X�̾�sҗ��cm��֯o'm�4Ʈ��f��y-pNyV�]�Gp�����ۂ5��U]<�U���<���A�r����*�V��~��K0�w,۝��Ĭ����	*A������Kdp���������Cp�`I	~�pV�Va�^ʹT�_t:sKrv0�y�xP���k�K4n벅�����ȣndG�tg߭D��o�_t�>��)�z�/�C �X(��Jϸ��$�;��}��7��R�R
�2��
�L*ns#�:�QB�yc�2K��o�N>Rх���c�o&����%>��S���y��C��Z��2��aԤ{<gb��"�@zJ��[ዒ�I��� ,C>�g�*��c������W�F��I��|���Rw@c��E-$��im�7�t�1�Cl3�v��@2<n�i��H`!Z��'�|8g�x��J=�n��2�qd���~y,Mޝy���M�'��gm�,�3�,��F�|o���.�"�95�O�'��l-���˿�g�+�%�G-�3�ߢ����?C��_�Mǧ[m��|�k���t[c��L{���{I3�DY���T������D�eH�V���H��`=�/J{]`Ⲩ�j�g-4?%/v �ʢ55�n� z�����<�0���g��2�ޟ4o�Tn���wq?��M9�	V���Z<^j��~�0A���Rͩ��m%��
�Zg��Q��I����2�\�6VtHQ'z�@.�9I��}/ɉ�����v�$Ү)�D�Y�6uU�#wr�cM��R�<Nez��������eѠ�>p'A�¯0�`?�ͼX^��x��-���[c�ӎ�GdqM���9�2ㆳ�� hAM�ʲk(`z��$I��9�j���!9 `��,�6$:�-�y�*5�z��Ų�����ons��)�7}��A)�9�QK�{,dޡq�h���i�"��{	x�铪���>���/�8N0�+A۟�m"CW�~p�:�a�l�PF^`By�LUN	,9�=d�sĠ���La��V����Z"�>��2��qJD��cB�R7�:�8���#��nV���t:�Nhr��Ma���f)9+�^��-P��ؙ3/�n���G���n��I%f+h.�x�����3�͎�� ϦZ�X�
�u<�qP��B�.~xE�$Y�����G�Hl���Kx�U�m�y	�6S�IL>��FW��O������AsAi�-���8�&# ����a��SJ��6��f�%��ϐO�ؚqƤ�:�c"���4f���Bu��.�(��e�7�g}׆|��T��]�O�k�ې���ow��IV#4z� ch-�2�{�@fA o�cM��ӡ��2J3wK(Wc��\��\%?�c!ŸUl�'����l�<�ۅ�b��C��.�iN�ﰾz*�g��u*�-�*�9D2��t�y��Lr1��TV\b��|�v�����ӊ�p��s�;i�\�]O�l�i�A��� �����!���!�������8r�W��#/�t�c����{-��������������A��!Gk0��Փ�t���f��qaVsQ�J������ܐv�x{	l�|���~~�,t��J��E7������C[.ӟJ�X�p�N^8����i_�����Z+�V|Y�D ��{&���ު��ۀ�P�%��)O𚼻D̂�,w��P㥎D$ܾ�h<���]�=&�ș�|Г�tOZ���R߿ T! I�PWS�u!A�톮O�R/�p�'�;ddq|G�C0�dgd��'v��u~i������\�� A�,R���{ۙ�m�����є}�,v*:i�1>^���و��S(6ߜ��ae�2>�i��°޲�\����t� �~A�Iw�2R��щ���u�����ɿ T��dOս�U��f���ܠ�n�Ṕo,<5 5��$q*N��7�:�s�+�L����evr�N�l/��U�}	V�1�Q�.�
�Phe���Z�ۿa�0,v�4Q��":�1E���փH��*&��s-	�Q�4��L��s��M}����æ��4Qf�%g�������p�G+��X�"���j�G	��>C]��۩Ɯc�0�A�]b�[���;�u�!�G��O:P��F��I�9��p/Z��'lޕ:��1V'�m�7�b��	L�a7�������2D)N�>��C��nɍ���zC��1dS �<�c�̝���=��])�a��L���ti�Nl�LlBr��yAlr������E�0W��/�Psq"J@KdI�#$N�
�>���,�?�J��ܠ~�e_�1�u/��ǧ��(R#�KO�3�:�&/+4'G�0s�1=;�Y��H2xZ��g�>�ҹ+:��[���y�Bu� fHNvkVRY]�S�e�0�5{�:0���$�ُ�^&L�k������`�qy��@�x����-�=�a/��Mǒ��(}�����%��o�D��y�#A� �6��|����eY7[05 �C0L��9I�E�K������fV#*^cHՑO�U��Pp�a ��1i�\�t�`��V�Y�֐A|������@�9�����ۅ�`�s�J �Wr��9K'��pp�꩸x�: �a�ݶ�$!�xBc��`g�eY�|-�=��o��F�H7�䟾dO�_L����w�X[fH��%��w9��$�~E셃�曣,�רV3S��]��6�?�~@��T��`#\�[������*� 9�kR֐��c��0W��5Y�,��1Eᣤ?�G9�67���B��6l{^����A�ȏ�0�:�@�
��o�w��D��;A��0��kbr�%��zUy�Ƹ)W�����3�k{NP��������_��1��T����<:Q���P�^ma�.H�#���'跈m�3�;����s"���O��}�2�/��L��z�f_�#K?����E�7
w����Qr.qx
��0��K��
��`�b�w������N�Xz��CXa����A���kE��B^���NaQ2���i;ik�
�o�QF/Q�_b=:6��0C�TY9����g��P@H�s���P� �����^Xs�Em+m`C�Vr�ŭ3��&=�����K�� @QĭT�b��ر�b/�ݽ�e�C��o�-�{O:`��h)�ƀO��s�ۆ� � Tx�$V-��3��L�j܁"U�".���r�`z�`V �p���LѬ>S\�5>��h�V����Ih
�ĥm�!�)�O��(�&0y�A)@_oJ�6A�����+w��!�����-t?he�,|&��d|:� %nGN#�9l�WsQ.��L�J�Ȃ� �`b(��ްĭ��|{�\�i�
iɽ����u�V�I��	������~���:>�b������_A�ε�����|�*U5�+@Z���L��*�/%��G�9%H�/Ӽ��Ae]��ח�\������̫�@rԮ�������QS�fїlO`:�',��EK�n�ڞ��!LDnٗO�����d���[�>r=8qp���X ��lf9)�DL/�S��р8{��8	Pd�&��Y��p7�?	b�Nk��&���טL�)��3���N������|ǯ�(G��k��A��2I��N�E!X����_�$(�AuI0e�f���]�B��r��5��5��<�S�΃�4$�~�d��=�/¿��w�L	ir7����S��+��w'�2��u������R
�(c
�٘���k�^H��k���_(�;�9�0"~)�,�Д�29�?��Ae{)��ja	���Nua���59�Uض���n ��@�����q��c���"��T�|�y��������G�yV5,�+��f��>�+c�:F�c�&-�����*'�/EL����3���O��e����a0�vﻱh���������u��
H�'��)VQ���=c�Eoh%�(2�������	ฝ��\'?�\+th�8K}�;,oA�㟎��e%`�FN9�M�Fe�q٥
/}��}(��"��;p� �6��oK-<��.�E���#��%3KF�2�<_lI�����D���`�b5�e�9Z@���Z�FD�(ڌ���v$fd�����櫫���<����o�iu �5�`	����7��m��o�i}����s�u��6�:e�d0�s��ө�O�*=��*��`�����8�ؒ�"ֵ]�y��n2_�^�%ˌw���߼3�a�Ϯ���+�Q�����&�T��i�Lx7�W�o�9�tw���)kׯ(���a��i��?\4
�ly�����'�vJ�x������&��N�*0��Ef����]jpi�S��+{9i���ؑ4�j��0vtk�/�x������ϲW��(;���Z�U�h��`�������}Ȉ�A4�U1�69�(&����5��#�L�)&�J;�A�����р*���i���
`ǺE�ą(y��_/*�`�3/�� ����1�WSeYH�UN�& ��54�_
s��ly�'Lc&P�E�JM|^�4�����Cp��n�2��[�� 	�F��Ծ�5��Kq�Q�Kn�y�F���&v	8����iZG�$W��]�+dPN��fC�����B̴�+�߷	����r6N^N�1'�&�Y-�%��h�?�8�!���_��M37��+���X໹�fh^�,��f),?�����B���������sL#Jj�2 E����@Ӆ[�C<p�K�Lb���Q�~\�W�W�0��0w����OQ@|��H7��b兘��@c�<ϟ�2<j�����F7_j��)�L�� n�%��dK�m�b��3��zČ�Ѣa�]�$�+>�{����Ҭ��6<|�H��sA����ѽ�să��s�H�
������S9�s��3���%32�G7&13�oł��O@S�}Lv�O3aG������p�8�:Jl.V��S#�!�M�+�#�^W���m�j�ZhF�̓fg	�&�n��_Ş��@�U�p͹�+��p��^@0YQj�E��a�L��5] �\��ڥ|~��L���2�0n'm�s}]����N/ԥĹH��@����R�ToTr;������i<��ɤY1�\z�I�}�5sx�FZ���^�N�`�wnFڌ8�ko�F���G���񄭇��>�#؏M��Ou4��=[��WA�Ѣ;)�����;*�L����1�=�K�`�秱�;ł]�僼a��!�H]��:��e�i��R#�{[9Z�g��N�!�Ms%Mg�aU,-n�h�"V��/��AK,i�aBm�&u4yn��p�qb�v^<yV�!� �Z+�q�,͘H!���rCbٳ%�'�$'�ʽ�c0��u(�06�B�� �)��g�.i9K�n���BͻB�bSy��м��;�9��R9`�n������q� ���	GK2]P H��ڗfɣ�o�	�_~r`,37���Hn!՘ϚN�3��w	k��6�тa�ꎑ�Q2mr;�
 AZ��d6�ܟݾ�W<�YnCv	447�Y�@��|��i&7��])p<�#>��)�����]t @� ��Ջbg��U�
�����s�����n���sP��+Xj��h���CCbx�v�O��Q�>F<�>��0�­M��s��m�7V}?���F_�Kr9ֆ�5A+w�	O�W=
���è?�ޑ$�T�{َ"���)i��Ξ�z��YkT����B��]H��/P�}-5� j74��)izի@Y �^9��熊	@���aJ�Y� ��G�XU�،����bu�����ᚆ+	�X)�v����/���� �+0+\�`�����[J�P��%���tg�V���8*�,ʣ��[c6��-D���6�L=w%�X1�|l�
�h�W?M+X��x]�.�*o�q_ŧf͐[lNE�Xo��}4���fo�}f��jc���ZY�?���΢֚���DW���:�0 �Zv���%5��gj|˛�`�i��E*�j�y#�ɨ�	�M��2�4vpY8Jk	I*���� �]V ��t�S �5���4L��c{VvĞ[����/�c�(ec��ފ�#˰��J�����N1w�����)���?��e�FH�c���l��*3[%�!��c1!/T�|s2f7���;NY'�]��?ų�(�M��҄���y2�@Y&ޟ:��)�T�@��'Дk��'�����nq#���ʞC�����1��n{���<��*,ɛ���ÈEQ��T��k��o��DyI0@s�O�@��y�L�,�;�F|��)O���ŕ$�f-��p��1������Ƚ�R|��X�r�d|��)���π�J�3#�$w�j��-��� ����1�Ah��O �<�ӟ�ST�����*߾gX5/�#�Z�R�=�o�-T��.���uF�ސ
"$���f��.qJe�������K��f��d~C]/�4fф��4���g>���9��P����o~�^eMT�-�� 9�X����!��W䌡��� c���i����d��箞��{W�47Y%X�>�ۧ�_v�ʇ��q����|H4�<4�2�cT��ܾ
��D��R�i��s�:?�z&��Fg��G@t+[c�<�]~�L��)�Q����(N���d��Cd2���CM^a+�Uw�2��wbᄦ	�7��k*Z;�+�5c6��?ދ)A2�`��}7Cbj�*MҔ��E1�c�D9�%�V��sı�)��� �/v&a�۴���e\zĨA��*+\!�H0n��K�b�j^���p.��~$'T�#d�_-i����7�p��,a��R�]���ꆽ�>�����!T��Y���۵��T4�,r1�Ie�BK���U@[�#)of��h/��.�ù��/i�u��H���a;I.\�4�ڙ��b_����7���i��7#�D4�GK;Nxv/2�k1����.r�*U�� ���y���g����Q�k�1�M{�_[Wm��pjfjy�v��El���R�w�1�)]PS��Ϥ`�� V��^L�];'˧�BM��)��� ��l�
�����ǒ�d�����V�IJ�뎤���x�{5P��4(LrG�f�u�
���ؘ�(�+9�tܙW���^]�7a�b�����|0B�(�;=Ev�'ҏ�ڶ�PL��N�(O?��/���^�ْ����: K*��yB-�s��]Ed���yk`A��O���fc�Z�{�"f�9%�3�-:���2��kwՓ"�1���^ZL� ���+�S�B�l?���0v�*lELĤ@U.�wZ"F� ���+�=,�+�gt*`�]�,��]0w����4�L*R�j"��_�x�#���OYK~��b��;;?���[x�?�؇�EHLrT����>;^e�[<o��A�yԆ�.�ͯ*DRAܰ�L���U�ͺ�i�l�r�H���%�U%P�xi�MLZ	yb^[S�W�!H�w��Ρ�z\s�]*ޏ�C:�D�'��4Xi�l�e��ǝ͏n�(����5�����6��h*N�N�VM�PpZ�ѧ�_-0�^���YB�+�C�#���	~ݫ�C�a�������@�9�,� F)�S���d�H���ֿ����'�+�/���h��Uxǣ�(k��P��܁�>��W�����>�R��b�IDͶZ�Z\B%k�j�h����.�U�;rX���	�v�_z�Hx�_w��
�N�Eu�	��)1"�-l��]�-'a�U���Vn����HR$f"�Y? b�H��&�t�T[?z�|r�vJ��k:��^LV9��TۋU�"K��+tR�X��m%�ð"����G:��������:$'�f���?��#�+x��S)_�%�f��ݦ���=���E�{�z�gRF��+�%�٬b���L3������!�5�����"h�1�?�|�{��_C{��\��^Wi��7zUF�����:�져��ق�Q�hk�����(�H"��c���j�">Vb=G���$�Jp"����e��
�HU�-]��HtC)_�}��]d����kz;t�|٦��1�u���e�1�Ň���1v�>փ('�K����w�HId<Ċ�f}.g'�mV����`�>Nc
��S�r���η&N�����O�:h�K		�hO��/��
ʭW��`��V�v�x�1{=@�l��xbɹ{�=�I6���'��&�w����"447OI� ��dò�л���ik�|�h`Q�kO&*��v=ͽﯻP�~��J�����Y�l�D����EI<^�F1o_�k�-��-��|�v��q��;y�Js�=y�\{6���'��u\��J3�	]-\cG�L9����k��ʀ�yE}��=��l���q��Ь�0i��55�4+��,��n~��;���W����@1V|-�SXZ�2�"�)�����bTaOC7�K�>W�5Er����p�q̠%�d �*#��#%�vr�B|]H��	x���AWi�sFivrr����F'���K�'@��v��õ���$F���)���=��-ۢ���z����=d����T��oK,;�e�N�� �	Е8�+ߛqY9U���Y�H�c�x2V:\����jg�p'-�}S�>E���e*�t�k���R�����L�Z��8i��#	t˴Wa������	�?�p��tSJ��kCw�E��,y퍏�6 *$Er�e���@e:��[h��e��7��"�0�l�	�L!��R�q��M��������K�����n��p��&fn���4�|f�.A�������KS*�.�%�7hS�O����N�]�T
VY�T�,v�J������8�_�q�C�m�諕��k eU�`���������g��y�`i������Q��9,���3�(��]�cp(����^��{��̫���Q՝a��"��n�8��ʄ� �p��wjV��-�2�W5����WQ�tw�;�A�Vdo1�\c��ћ�^@x�!�b�t��.Iz�NEѨ%��5��	!��	��9�ZM�PٗϤW]�YU$����ݨȤū:r�<��%8�C����ԳW5'���G��y���$Ǚ�.��2H����V�'�X�Y�rI9���^�[�A�	�zC�d���i�<�ME�8!��Jr��1������?�RI�OIW�|�G�T�9y�0�BPW��,�qYo���I\-�_��CH��E�"^O�0]p���?�xoYR�� #���ȶ�2�zJ�mgG����zd�U����1�Ľ�D��9ۜ�0����|?�b�U{H�X�}�o�M�;Ӏ�.��۾�Y_;ƛ\u���6�'��a��h����H��v㨎b-�*��z���f�*��u�J��Ɏ�~�_�t�"?�:�vDD��Op(n*��~bA3!�H�HNI�;�sI�$?hC��������9{�����E�pa�{���E�zj̓j䮩�?-�܎���y���wl�&Y�v唎k�;9&Q�:�V��w?����7�9W3Hՠݬl��V�Ϊ��n'�P>�J 3tv�+�N�Q�R�&�
�����ql�k��+e�6FB��ɂ�!h�ػF�Lus`YQI�2E�%h�n�.�Q�+��Q�B$G�ޔ�ȫ��A��IT�ܞ�y��������^w���eR��n�p&��w95o�ou��(���^�	Isoc��GrQ���܃g.�x�7f��P�U��Gɓx�N�/#�v��=J?��$v!kv�O[I�zJ�E�k��h2�� _��PwBM���
����9BwTx�xЀc�O�E�J��l��~�dr^���pcF�
�ip|��C�ִ�'F�]D��l�o5�p�0����U���t�g�^V;Eה(����tl���e�.�ŵ��^V���y��f�I�����C�˃'�(�A�ƌ�ņ�,V<�Dp1�oaON�����R3�8`������2	eg����qux1�H��	��t��F)wΩ��?����_M���C��m���-	|��	�������2��������[֐ߧ���&OUSR���>��<�æ�z��� �{=\ )[.���X�^,�G|�]N��1jF8���m>�%���AO(�!,i���W��M%�Ӡh�L�<���� T����s]5� ��)� K�P����}&l�6�B��nÓ��1ug���Jw��?�+�J}��Cǈ)t�R���9DN+&0�|��A�d�an���@������6�Y���L̬�:��jY��	-ϔ�|��9gBr���Ӡ�_	v%�k���9�	�1d��,S���:R�@�]w�)
����p�����e��b&ax^9	�P+{���\��-��ZwtVjm�o��b�9�]�(Ƽk����'p@ϳh0�|+��K�P�$��qȊ7��>G:������2e���۫P.�nr�w�t}�&��c�#r�:{~zu8��A��k��@���6.jBx5q�u$vp�R	b�kN>�7zQ�ȲPoP����f���f�W7�}�2P�_�:x�Ͱ�#�����˙_�Ś����1�Y�tt��Dy:�E�$l��5��̰����f�@"��yH�2�䠉ղ5�D��%���%�\�gv?w��I�˱�,���,����t�
��U>�v�ǣ�t$��#"�R����S���|��J�r?��p������~��s1��s�r�-ǦV��R�Y�L��~��[wV����
�
�; �����^��'��;���g���l�)^�l��>��c $�s�0ߵ�A�4(wy���3����6j4�	k���S���%Y��Qֿ���RA�M��{��44$pb��yB{>��}��9�������z�æ����DP�]�.Z�G�8���=��U����D/�lP%�w��ďԝ$׍)*5�&
_�T�*݂&�َ�E�*�y WRX//�}��9��g�?:D�G�v�S���kd�KGꢮCFÀe��Yz��һ:�7��9��Ž�+�3m��N)�ɤ��P���Yi�.��Ƀ���	؜N���1�Q�n�c�_�1�n�^���m��L�"��ka�Ȝ6�}0�B�U�p��O����ŋ־���k=�f��Ý2�V���������81��s�	�q	��5K�H
i�2_FZ�f��^ʙ�p�YvzQp������I�Da���Jw4&�4hi���-���V�с�N�n9���4�*\���C#]�$cTMR�������n�L��P(ޯ���Ψ�=}�c���+ޞ�3�Ԏ�.���5o~�X�>�[zTغ���a ������U-�m��i��X����;�c�Z��-�T����m0p.��� AA%t�ZkXQ��J#�R�V'1VقmzX� l� f��VT�pX��uy��-�`��m���W%w�~�.{%*�Q}+�-�Gڝ#
�.�ve��ǯ�]��+��6��_�W�����㫸��G���T㯑����p>:W?��n�#���8�bf;�o^�����UVDp�N��w�5�iĻc�)�c��,05�-b���o(ż;��.��x2������y�K�@���x��@eSA���$<�
{�q�p��By)���#�j]���w=vp�ݭ��u��T�t��%ny0�5���>w�?}����eʔ�gu�Y��?��^*;3^W��82�3$j������A� ~���C��3�t((�p"dc��:�;:����<S�<6�#Ԃ!�z^�	�Kc"��U��(��c��R1~7k�v��E�tO�VE1 e���G��L�=�������n?2���X��Ӷ��~��THǰ�]u�3l�I��HA�@��X	�O4�4��PP����D��]���~�Q1Ar��7z�`��7���!��(�ҝ�THA�P?i�t����H�� �sR浢֪T�g۹z��3�=o,˞�}�'������ )T�VCT��E��6�>o>��%1Wam^�vƥ�DQNI�Qa�Pf"���̍�#���8xї��瞫�T�7��mV��q���w��(�v!z�R�ѝnJZ�Lh�|N�-��0�i_8k��d�x��&F��dڜUh�`����^\��k\a=1Q��A��T_>�Nf���Vi�1�	�[(�97U�d_�	##��, �%,{�E���v5m�F�����ZI�p�4��F�m2l�>�L�b��z��/S����0��s�i�*�/�К�[b������/R��D���[�SW-�ir��Lw!�O����bCB�_7�c��I�nA0j^8HT�}�����!��`���`����x�zh��jy�:���.��=��a)�˫.e�#�nC`f�z��ܖ�H�F"M�@�aY�ϺK<��i�0<-��m��;>-��%CXOY	��>ˆvYe �!�F*��Ə�'�cS�zB:�uA�|������0= �D�h�M��>-��T*��OIU{�(O	���yj�A����j[FY����������j�'ٺ42d����=�m�zS�Ȧ,9Q*��%%~,�J�C�^>4s�c���_[��7�.g����E:���
� �2uF�)"�~;��y4��G��V�4��=ј��!��B(�M��L���������Ɣk��NI�ȍEF'�P�(�N%�B����/�����%���	Xݥ�υ}���G�n�ƾ��_��qa�="R9���������q�G�ك�Km$` a��C���%=�XvD=an��f����Ⱦk��h�aϊ]�V�Dl�^t��i:A�2.��M��*^$ih*XY|�Rl�LT�,����m��4Ë�yS��a4Jd�k�!%�7���?���7��(�SJ��gb��g[����Z��/-jp��ǯn��ae�ɸ Y[1�,�uZb�2�({�f���4�T{���2l�0�}��'*��ۗ���,�t��e��a��38���&�N}@�eo�����I�&��c;[C.i}�r��Ʌ���I�Z+��*AM�AL�V��hK9k��[�����]j�#����R�X}���t4 �VQ��]6�q�~���s`j�
�N#,��V'�0���
]�D���&\U�?���ہ���
�,�=�=]�e7�ǌ� ��[$Ӝ��q��qT��c�훮*t?9�}��I�-L:HA���[y�m	�x�e��ؠQ�ǀ���ՙrQj:3�=��;8(�ho�c=s��Xd2]�ԅ�������+�҂Feu+�ء��E�i���h��x<��X!ʞ�*�ҽA
���"y��R2����������x�+����{(��׍�X��k��=�C�8Po��բ�׀������a��D���u����ĳ�q�0�OOq����
`���Ł��A&|�c�OZ0�"�&����.�j��¼�V sY��[�"��@)&/�ن�k�ʕI����)��'�L����An� VT�ޡ���ݫ+'Q�_��.���n���J�P�Q8��6�����.���=P(
�F@��I����\`��P2bx��h~ܓ�A���Q��'�p��2"�l��(���I\�)!ܕ
؉`�-8�w��ln��9S��_]��*\B��>���IkI4uF/��.�8�vu��1�Ѣ�h������]��P,�Y�
ċP"h�eI7��÷��Yh�5��#t�E�=SC H�DZ��:��TBb���'%�n,w�J��1�{�&���ꋳˣ�P�X�*�iiEQ־�
���y�ݤv��]v�-��	d��]���<b��!NQ��J�۷���C���|��.C�W����.���Q4ƅ����]*��眇�W�Ki!��^toKS���̊)�ur��E['(���D�țA�|с��(�O\��)��U��-�yھS�h.�Zй8���4'v*�FV��>r�_Aa����E��cBә�[v.�2{����j��,T��&�L����������O���Z-��w�RK����=���@��?����Pjk��.��OBcߣ��"Ȩ�R
����0�͆?(�6Nl�=���Z��E�3��w/b��EK7.�,�к�R�ԯ�HL�yD�Q]$�a7�n�=y`��I��f
T4z>���Y͇Q�{6#SS�W��w�S� ��9�:�
9��%�q���uiG�	�O��F
 ]�<+͚�}�I�,��Xu�Z�1�`�-���J��0<\7lY�bF���||(l�����'��0|�����7A`T?�"$y���x�6�;%�H/43�z3�mr���C����j>�34�ߚ�E]�[StÐ��O�^��D���7PC��=����=p�:ޕd�-!�h���ŉ!\�]���b��@jp�cU�3�6��l,�Y�T��Wn{Wl�J�{��m.К8���+ײ$am����霢e ��<�Q�X��J�j֯S�+��"D�B��\i��P�@��._��+�����Yڹ����(�ux5'�p�(B���9�o���'߼
�M�:xߥ��NM1��ri���j7BW�8��\L9[���+����i+B��<�ܸs��Y��&8�]ڥ��P�d�@�+[l,}��-�_$y+·�g��z�V�l>�V���Kߞ|n�����m}��&
H���{UȦ��%g��㓔�'R�5���:�-��#� �v���M��T�$�v?Q�3es��?z����$��@�ejHFCs8/�����[Q�<Es3/��}����CyI�9L>�l.�;�NX䛕W��~�H�텷�hCھ(@N�ۜ�?�j���܊������<���q���J�|qSE�`��p{x{�f�Ҁ��t0$���t>.�i��j��h�`V/������_K�@��Lj�OI&�3�_�Wֿ0ƴ�2棒�ZF���f��αâ<���e����N������sg��Y�="���n�~��/k�G�30��.�
L���"~��I�M��ׄ�7�C5���YZ��=���Y�7(� �'�(!�J����L<�`M~�a|��0��M��Y�Y�Av{dĠxóq�7�񰬺����'�$˺F����	/v�_v�9�͙�OJ���RȄ��Į�X=�_���T�:������U��5)��ĎI p.yu�qڃ���UҐfy�wr��U�/�H7�Qi�G-2j���:x�"%�T�9��x�F�O������E��h�0X�v�0����b	o���ga�_*�H��,���#Bי����l�����<�s�l/�"�Z��s8����(��fy�{뎲q�z������a�0�F4�L�����$�K�u�Ve�*�֦���@�|yX��˧���C�v�	�&b� ��Ð-�A��1��!�c�������%��?[��a�.@G2x.HsA�п�/"��GU�`._���>�zr,9+pu^����r�6?�&r���Jgx�;�,ڔ#���vT*�>�Bjg8)[��a������D?��⣻}r�(0���i^E~J��G`\lv񄀥ء���z;I�H0l=Ȣ�r0��9F$�w�k��w�Ҍ�c5y��<�k?±[6`�m��)��m�1L1�����䭨P�	���@��¡��e�mC2��u�`���^��>�?�R)^�^�F{Bc;R��dp&�%�ar!Ly�%�L����A5��;r��r�kH�20m6K��[fA���p`�/%���T�i��ô	����ޖ�By��{��2��h�u���c��	��&'μ`�(i��K���,��Ϲ��I����E��pTW� ��Lc3d��3�S�ߜg+%��G���b���^��c��`p牋\3����%�=-��'T�����:�c�Ȩ�~�̛SG��s���CR�$����h���G&Ր��-�b$�w�E�h���t���X;b�y�J�
| � ��_
�¢��␓�<sv�E�k��{
�'�N>��]Q�^���}D�
n������a�P�,�k
:�-�2�5��*�N�j�:Q�5��]5OV�X<�|��V��a��	�i�d|�rn�hW��M4r��Z�2��7LJn�-ُe�xNL4��/+�Z�H���������|���1d��O.����B�
=9�]�\��T�)��Y�x�M�JQ"�৥cN;�7Ʀ�<6�iV�e�2�T���P�G�Cg|#��D��!?mVj�<*�燚��[t�\�r����P �g�+qH$�iX��܁c�L��9]8�짯��Kn���}&ʘ0	����V��s�o��ځ�����:��Bk��Z�j����h��r@���̱�^Dl�����C��k��X�e5���D�'��s*�5�}�H�m�5;�c~So�E��S!n��������qAc��5T�Q��V�����^P�������a9�cZ�N0�l��d>$�/�sO�������xK&����������m2�r ����z7�A�����b���m�H<�15��A�>�e~=��ȏr��f�(>��b�Qw��p�ckK�0�,p�ob��}�.�⡠EH�ۣL�M2�A[��v��������)�`k5����*���"�8XB���>\F��O*%
��"�wL�!g`M,o�ý��Wg�P�ӮÍ���@M�b[[CF�z7��#��v��i'}�ދi�Ϳ3s�Z#P,𜠀	b���:^!����r�6-'������9᪽ӌU�2�,��8W��L�s��_���#q��EC(��=�P�p�F'�e�R�qK`p�[R9��q���A�q2��5B����3��b��Ѣu��t;�+4<0��C&堑���CeX/��y[���%���Z��-�\Aٚ�]%���2��r��]G�C����t��мo�2u-��?�t��u-t=[�gj�fK�~ɯz\���˱��<�!%�ߓ����|�}�o
�kr�|]9�H����Ɯ<g6"�%�TI8c7H�2+�q?� �gL1���eIeɷ��.3���TMP�Ջ�co;q�.��>��B �r%O�!�.�1��!�^��N����x��w7�ƽ$^5z\.ڜ�Ϩ�|җߧ}ʶ�l7Oy/yy�/m�4Hu=��>!�=1�J�k/`[�&f�h��RE�F/L��(�-t��撕�>��Cps1��S�&�;pM���!���q)L|(���0��;5��n:��l���rb�
����	|r](f�P�ٛY��mL�!̥+��рg�L�,*�V[�@\a@���=�����&P�βWƔ������r~j���Ť���W��ۮ��?ٓnr���'����w 0�[.WX'M5�w+y�8C�-�lճ�]eTVCk���)�ݭ,�K�I� +	�٣�sҘY�vQ�<8S�WJ�I���n�&T�����	�6�-���T�N���������ͤ��Ş,��c`S��h�7�� �|p�ҙk�0y�j�ow�r�F�\�X�?�)_��.��h�B�DW�B�s������|��<[G�c�q&:�@"Y�J���@#���s������M&�A�Vz�I`���}|���u�/��E+�]�<��.�Oo{v�lȹ��I�O��ӷ{�-�l�dM:���>tk�Ƥ��
�'����0�z�|�f���tx������e��@��a��Èm�ͦ�Ds��)UX��f ����WL�%��TN#�����(�����X�I�g�O�:�� �W�w[�rA��l�$_!�@��"_��'������%�G$3�h��w4�x�����A�8.�����k^�'��=��0� �L》^S@��Z_b�~��&���9'�Q+��v�C;:����r�o��!��7n�,�X��EsZ�ך`��]�"�E�|d��*ᇹ+�I�n��߾�|>�#�g��1�#��ؙ��RL*�z��v@��CM�HD��u̢$�!-G�AK��t#�����g���Ϥ�J��Ѳ����,W*(a}�Hx�ގ�=Ҙ�,�NgB��n�$��fN��­|٦�U��� es��\���W��5��pe�,�lϽ���О��'�:�1�:zoӻ�&�=�����
��N��4/���^�L�Y؈�Z%�g̎����br��`�������� �Q��pO;��BY��>z%������/�-@WȋUzq�6��1���t�����Qh:�Oܬ�ܚq��:���S}���5�?�����V��:�hy��Д�; ��<��g���$����od,d+�1�Ÿ�5�x�,yfG2�v�b� ����x�]�zIX�M3*KH�!�<9��|a�C�����q�Eo�o�}Cm��_��k玸o}4��hhH�y��5EޠЦ6u����������]M���7�-{�ͮ��{|���~���Z��X�C��}�<+i_�½��՜h'�<!�`�Zz�����o	�<��)�śf#��	X13B�o�b���d�is��znlJ����Dh� 5�l���o�8
ww��Fż���f�H���D�gp����5��0oH��l�����U'4�Y�^l�=���Y��Ij����faS6@�7�N��(dQD�Wm �8:�~��_F���o�]�f�0�M@	����ɅH>6�_ڐ_sDh�a�ƀ`r9��l�Y��������������4r\K��2�A
�Q���9u���v�o����p��7�c\�B��o+�FW�s0�V���{�(��n�����v�K�S��F@�l��������*��O뙔��$�*�YF*���`���\)��Wn�����fY녒lQ�S\60�������J{j'Q��� gOo+�y�w���~h0���SY>�LY�}�	��T���2���4��w#)����ԥ�O�K�Kk�J���I>L�;�B+󳬵�cT7��X�J��o�	�qqx�R/������c���$K��d��ԕŌ����p���V!����W�H�M^:T�N���ִ�+pC���H�25��B3]���i��.�Iu[,����u�9T��Q#بT����m�
��d~����:�՗�WuY�M�Ipd���6�2hnZi�*>�S�i���7Z?iǺ�=L���S���H�Z�$XH��!y�$rUح��E�xlf_C�qj�̐`���i�V���~V����@�c��yгZ-g��b��?�2��߮,�Ut��D.���U{X�Ju�1!z�io�9�X8yE+C_�k�h�,�r���	U&���?�w��Tx�n
cT۠s nU�n��]C9狭p����$����F�-4H,�7�B2����YւN��`)44�-K�#d�F�c�7�0:���&��v<��6��(P��e]�2h���^V�N�IЁ���0G�`�é�'�A˩��<��'�tq-)O�~���� u�b$��N>����x`!����0x)�����pw�ȿW�H$��C>�q�X�:.���Șo��C����d5e��{����1��Pu��}����+j3~�hI��=A�Q�$߰��4�;?�3棳��Gs����]�(�7tbڎ��Z����w?LwX$Ҭ��1P�/��]�t��)j/���ukf#�d-���xgX5IY�%h�U	kє�&��N�'��6J�g�{�;�;���%�����/��xƯB�N8���R�w�X٭?��TUd8�(����-K9K�aƍ��nܕ�qUI�0՘�r���-�a���*�wvL�ܥ�A.?�ܾ@yP����ΐ��Zt��b�	$�+~-9�j\`=Ƀ����qF�5UF�꽔8T�� k'��S��u����p��$Ҩ~����0G��s��W���Vv�>U�Eņ�J�}�lj�S�^�q�ec0�[i�
���rTae�FH�[t۝U����z��i��(��.����L��îZ��5x��/C	@y��1��R�mpm�J�V����RC�|;���j�����g)%:�dp.K	�~V�*�_
U�C'(�N�����6]6dOf��Hw�^�8��Y��%Jۓ�GN��颮���̵���bW	`�Ǽ:{�tɝ+����I޼�g�>�p���P׌�!��/9;�E���G5��7��A�������������|V즒�/?���\�U-���+_5O���U��T�"6�k�����-<ِN�T:�����;\��X��)�篜X����-�_��<F; ���i8d�T�?�RQE:�>yj|ݎ�|8:z��3:rk��Iµm�˳@u	J]�hDH7b�u��~��jD&���y���"��B�E�@*�VtB��x�P��[�iX��"��a�_i]\�8��5�`0j��" ���l�r�Eg��9����i���H|���.P�*�un�y
]n���q1(�S���	I��U��ir���8A���B��ݺ`Я:��$��xZ��3�s�p�Z�4E	��"���fmc(dBy�I�u_�sOܝa#��Պ�rUm�&�"�`��5�A�B!�.�/��~�QNNu�$����=ȁ"����u�q^�����~kj�y�BT^�S�'��V�J\�g4u�O�PD��9��f�}	e�,xHC��h�IH#q���ʁP�����S���&���4z�{HQS$������J��͟�3��mnP��R�W��`���\F����qb�YN�M��.9�%=��-�O���\(k	�{']P2�Vh�1	F��ܽw��hѲRF��g��[�
���2�0�1��ն7�����=\����ժT�;�!�3j��l#��f�f�����&цk&���6���6��(0b҇��8�3x)Sљ��0(�"��휚�BnkgZ3P
Jcy���55
�sR���� P�-4߈H,�C�� ���F0��	�)e� %�<{F�8�qP��Sd[[����o���]ȄhkхF���&���XT[T�7kw@q�0���ʹ�5��^�'ԙR���5�8��sB�)���lc$��9�b�AF��M���vᾨ"1^���S)(���W�El��ъB�����#��)LӾ�!w��w�h�e��M�Ш���Zu<�U��0��R���OV�I������G�E����5��5��a,|�;X�����>����p�`{lR�éG���F'#U?:�bv����36�j����Jqb��n����� =�Y)yb�c�g��l�[��&�@V�7���xR���s3&�&����L�"4���UQ��]�ݺ����U��Z�Ս*7o�;O�,{w;�n#�qU���|:�vY�ՖK
C�ulz�$�_{�FGdL��!��՘$���.qu�E3��
�b��ͼXއU3t�cZ&/�6osVA�������+���à��¿DX�Eo_ƠVo�[�g��
�
�DyI�1/=<��;u��!v�F�T|k:��mO�P���Vf���j0)��i��5����`�\&k){s}΀�$NN�~�2��M%)w]�.2��˘w��"a�M����&�*;�\H\�E7���M����=��c�&�5���u!S�]��il�bHn��)�)��(
b���
�#�'�3�c����! P
6�+�^�
�хؒ�UY�a��[},�(v�$:ًB�����b�������Q�<�z���U�HB
���
A��	Τ%��`�,)�'H»�f-b�s��3vD;����n�7�d��2/x��m�\�
}���M�G9��)������i�
iG%�{ ���b�z�F*NP�<;��*=�S������dt q���kưƖ=��D&R���[�$ =yohQ��͢��R"���1��愢��Ń;I���q�|��R�X=��W ���,�c-K8/��wQ��.βd=�	_;{�=��^�ȳ�/�Lfb�\vt����/%fA*�#�����d`�`շ?P�rQ}h�^�܍E+!�H�Lܼ�v��1�b ˕��	��H�����oU�K(�O�������Tҥ�yi�gaP���z�.O��KPt� Y�]2\e-,�Εql�YE���OP�p�I� 8v
���
*�4#���\�����bmm�p�Qn�X��v;�D���d�	�i�I��5�ݧ�u?n����F�0�:.y��Z��Vſb�{;��>��y�8 ��H\2y7��]��P��U���Оm����Q�aVJ��<�	�Dg��~�mR�ǱY��H��@��������x�xT
R�"0H:�o"��d�W�S����˴jʘ]̆��m 㯞6�+h�n��
�|�gh�a%� G�l��Q�;�B�Pqt� c�=���N����'5��ѕt���.�3��O9�I#��FA�u�H�f�b&�!��!c�HM��q�5ђ�$��.�����fnB���`x�6�62Yf��qZ��i���=+���?�er��*�7
l5r�)�oV�87΅�UEO�/�
N^�5������趡�>0j�~	m^��ͫ���ȪH�N�⃈1#����ʂ8����mYdK��.�r�����l����Ծ�ke���
�������-�<�
�E,RDPd0�稍&hq�'���g�c�����kiZТ6�J�5��/JQ������uh8IX8)xMê�2��kn�%+��[���ɫ��%;�I� ��C����5i��VRnrLl+��|�N�/	;�*L�ńJ��!T��\��I����Ea	�����NN��|H���I��r��+kD�N�o:� ���#0͞�.��5��ğ@Q�d��f��5j6b:�3\���B�����;�B�{e,���@�E��S;Dv�_<�ȟ��H�`�`��3[/����������6�+��¢�ٹ�}�n�9
qf<qK4_?����h�����!��Z1TL���רM���W[?����	�,P%�2�h���TA�D�bK1"g�+ק��筱i�țU�&���Q_�s��Ce�~R��C�Y�@���<�w=4E'/n�7$��a�k��^����紆хq�0>To�q��e1" ",�hd=XX��:t0Ę(�׫f+����Ӎ"�����[���L�j�b����?s��'hL�Qj�5@X�ْ`L4O�O@BA5�A���Ib��*�Ɩ�*`�L�1��bA��&������w
wGf�c�W:��0�"NV\�z�atL��ܛ��w����@���x&�_*�*<E��q���ذq�*1���'��Sf���k���k
*$�Jт��@�����J=k��cw@��}ݽo�V�N���I��j�C�>�&�碌�l���β��������ϴI\�]=D�L�t��}@�T'�y4c�\Y�����K����`c�	�1��{���D�&=�����kҼ�6}�E��*����{��ğfl�<!'pb�s��ƄF��ۥ^y��|..`���ܦ�����"�#����@6��%�� :K��N����4��Qf���t"~f���"ᝧ�-��O�k��oV���rO�2�|MO����P��9'D:,�qޫ�j-�4I�Fˎ��q��ہő���tcЗBO!f�B"�x6�y��H��fu�O1/YQ�J�e�b�8������Ĕ�7��^�,�JQȅū�]=����p'W�^׻�q�gjVN7�δ�Rd��H�`��좞#�$����LK�[����M�/��jV�$.�e��-�4k���P�I��O��/@Z�+3�6�ꖬ�Xѝli#�d�|4w�J=Gx�p�_x�����K# !�G�����71�B>�dt�"����<6X�/$��j�[h���F�9�(�h��K�y��L��J� �$� nk<?���xC��>����Ux��u�����;v����W��rG�|@ j�SB��@gش��%y}P��u+�@K�!9��*��+�7�	5�1*��������p=IC<�:�ء���* ���f�<�GCvC�j����H�K�%�/R�M�@�������m0O �U�b�0Mw�(q���:����S�����|���2;�>�`Wk�`tP�b�~S#��0.��~�*�!%h���M�ʁ΀2�����{�FXP��yB|T�P��;�M2�\���g�\>}�����/=��/aݑ+'Ĉ:=��?�{��T7��������>��"��G,�yL����{���s�F%a���{D.���k�cuw��a�]X�s��A_�j��F&W$H�x\�Ih�g������*U n]���:�	�n�e_kmA��@�{U�g0h��3��v�^.���H�&�ƖF�NY��D�P�����Jĸ�3o�����qf��G�&��Ƹw��d2X�Z�����Zr����v卾��	��08D�:%Z�)��X�A�P8U�[$K�O;��A�������~����1PX�i�1��B_�Ѹ֟ܜ^��1�`�H�I�j_�?s����p�w�Ӎ ��ÜQ;��+��*�L뒪ZG�f]}����(/�ē*�]+���#uje:Θ� ^Kz�,���،�v��g�ψ��7��OL��;fѿ�=��S��Ȩ�~_*=���Q)�ڰi!G��ĉ�
��#ֆ���t
`�!C�~���[�%�,	`��N�IСR��UR
Y�1wÙ�ׯ-7��[EMN	7@IM�#���9_��.�a��� &��ł��jH�qo���`Cf�[�u�7��\�`�!Sq9ڸ6��B��e�C�'r�A>}�^)����O�p�\�Uh���$?����3N����-�r:��w�P�+�@*�-���8'Z�7�q;��_�`���{�2g�x��ި�J2���j`r1?Qj&�Ma�H��)��q��x.�6fUQ�������TsN���g�B4@�x��㦝	R��D5�7��e��̰�"H����~�P���w�^�z�n_(�wƔq}�r
a�����J��+�O�l-e�(6����qr�%>|�]]e��g,�ZO\�!"����1��l�gG�"�K|��d�����gʶ��rS�esY^N(��(�xH�@A�f���� �0<BuЏ7�PR��3����E���#�Ȍ_j2�_o�|����b��اwg�!��qT�8���g�mV�������C�H����Ȥn�<��]#�R���6�088��\�NMf�H�e5�}���0�����(�Şo�!&�d��Jh+O��'H���ݓ��U���x���w�|�������9&�y��Jї�g�)�]�������H$PB�@!Y~!�������5�߈G��U��띓<��wyG6X/"ĺ��2�#wy@p�Z̭��͇�E��z�lbl� ��J���R����Q��X��G4�<�g@t��b=�W��D�(���Z�t9*\�%�h��J�|�+|0Y?�r�fE�j�K�P58\w�AH���r>�
��1$W��A�1�	_3\\�(�ˎ �u��*B���E�Ѭ���S�v��H73�g��	`]+A��s������R��<0d38�n�����}�-Ȧ½C���U�ӝ|�^0��ih\��א�.[!Pp�Lw�[h�F�z�S5h^�QOj(�'sQ��e��g/w@3*qIHHp3�҂�&i��V6R�%B
4��CT>�߁��Jښp3�i7���&����3�rG �>�X��."l�@�x{3;7mt�yVխ�,�{gM��8����Ò7q��A��d���ˎZ����o�K�3���t�P�a1ƴ����J�Mu��8x�x9���zO�(�\�E/��������=A畫�;T�T;��n�W��MU;a�u)��%�����	��;{��>��٪f��mz�13.4z2<.h�\%�]6�����J�(�{��U�����D>�-$_�)�	y8�xb�j�_�}� �)�m����vT#�|�<븥]a�_�C��ݙYT��y`}	2�=�D2�0���Q=�j��6��(L���{V��R�"9[|�� 	�Z@Y�w���.�.����
%���2d����@Yʱ�HKU���/`:)��yB����
�ob�7���p-��A��PS<n�'qr�ui��(�m�\Yc?J�wӡAGL�n-,����rL@~��#��x�}�W�����ZXi������\��fGhя\�e�g�����jz��݁�&C%*��&ާuXZ�y�rr�VW=�gY�B��Bv��G����
 ���񘊬l�
J'�9.w��?��ԻS)�O�0!�w��`�6уݜ[���RJ�j���'�#N�L��tL�?!�z�ٿ �hU�XIJ'�p�����+���+yO�h������bγ�`�_\Q!.ZP}��˾��쟏�T5r���e�	�*l���iq�l��bўT���U���O�N���Od�wZW�Nn�O������@1����8ܚ9�z�i�$�]��}Td\�� ���a�l|:C�C	X��\������e�`���#��/e�:���G�V.�jlև�.{�vL�ӌLڟ�6k���ƶgj�Bt�m�*�d�c��[����s���x#[��K����ƣ������l��ZM��q~$:�5�.�c��׶nP��� �Y�1f^�X9�S_��L���6��Aj�1���YX�#?ԑ��r!��*�+o�(E��?6�/�P �2�w,��9�i%��d�[2s�R�:�6A|Σ6w	��K�[�5vMYPx��,�]ca�*����KI(A���}>�-�"���A\��U+~@b
Ֆ?ǿ���TX�Ա�2DT��
�D�ߌ�"5ck'|f�{"�I$��i0��-�HL���R�/LU��!��m�Mw�A_?C��:�]g����6B�8�����Ƙ�?��
`f��f�ԣx}Tqv<�b[��t����W�W#�Mi��Yt�:z�B�`?��xn�Y�=F�*l5:8J)���{1j�ᚴV�O*��<�AX@U�%W�u��
��_}���j�t�L�j,�m�?澒�MY�8r�ʠF�{�kӣ8��:�3;
��C����ϫ��>��qQ�lKu}fm]8<��6I�-��>7�~�,�8�ep�*�͔N��?+�����ڋ�e���Z���ʕ���W�� ��̵�5��t�a�,pWZ��@�!��,)M;�p�`���	3Ҷ�H3f_2q�bz�y?�W��t����_�����/x�6@{�g�2J��?Y�~r���ӨE76:��>D�alSU���/^��F�U��l>o*B� o��ݓ����|X	�dl|J��R��Z�l����aD=��K���DFT?ĵllM"���׆q')Ǜ��-�]阭2��������ڒIf��$��c ��.�ӧ
��������)����d�K.z&ķ	5h�r�j����B���[ ���Pǂ�����o��	�hz�:�4�x�����Cfȹ�/p>��?�T��������e���ǰ�_��3߃��$y�Ɏ�n�%�tgG^����]f�.�KA��ج���X"rݯ9����[?Տ\>�RpN4���R3���#����I�-��%�;�',��S����Q'"�5���\|Ow�@��(bb��@�`TJ�ȠU�}Dj
e]�����Jeةާ��� �������ίW-po��V$�Tw�z.���a{�T;~��>�Avߕ0w��W��13a &�RW���q���_
���G����Z"������WE�4U��s�	����E��	��{�	g��o��c���B'��F�@��a��В�g��.QBTe�ǂ�(�XP���U����q^U���_�=����2lZ��������ɿ.�D3�{a��)�u��)�Y8s�X�)��Y��nu�@��5��R��-�⺫&�V��3�3���*\�C�6� K�(�7����/IM/�%���Q��.��W:jjBv�����bǘW���	��7D��lt��2����,%�
�]�
�)HdO`�;������$v��b�_N�IN'�#���ER EC��:!�P�⩭���sv1Θ_ZB��Y�O���Sj������2�U=g����^�n�[#�%�P��BR�	��99b�%���4@Q�����*�+���ip%_�}����\���	��}Ŭ���������)7�r�'�:ZM��������]A|�ѵ� �Z\��9wlE�.���P˰������ �[]� ��j�}n����p���� �(�V{-�pl�dv���}G+��U������#,��S>��)��̺���j�)x|&�y!DbJ[���{(r
�U^��%؉��I@����}���ě�z�x����7;�xDv�}[�a��w�}�����"���l�K,�s��l����4<�/�
Ī�<9���d�_�U+���ů������9��訉�������~��8�H�_��LW���JkN�s�Hֆ+Js�<A������ �����{Q�M��H/�6�	t\٪X8nq��:J�a��H�t��Gr9� ��V
��ڄ�&�D�wW�Q�i����9�!ޏ��4����,�����G�H�K�k`x맱j-��\���z��ZB����iOl&�K*�}n�i��?��Sr`�b@��-��p�~�}�lGǿ�Zү�5^���#�g!F�R��av��<HN�C�\Q���ﰆ�ϣ�H�HL D�F�|$�Ǌ�C?��Pd�Y5@bZ�R�ȅ���t1���vF�,���:�M��W���ٷ��&�g����G�����&O)9ێ)Ž
�V/c:#��6��r@O\"�0`�*!<i�s��;�d�g���Rg�6z�VK������x���7��������B�TK�	�?���A�WL ,�BP�Ta0#��p(n�j�~�9���OT���V�?=��@���s�.O�)���C��D�n�.I^*U�r�����(�rgp�"���[4Ü*�{�pȑ��5�F��>�ޕD��me��\�*�՚8m�⚘����p��Mx7��R'����Gau���i�'"i����� L'����&�J��:.)���!*�o�O�cu���_���?5#[K�+�/�NXF<�??!����P��[œ�BzKu��?���L�*@Q<16}�������h@�gv����T�B0����@C�`�$�wwr�p ���� �g1/��=\���1�LQF׃�wz��b�,���Z�Z���%� ���nXjv+>�j�I��wWO�<�~���Á~�ji%e�g�L�0aL�#���%����>BVU�/�8���t<U�WL�E�����f�#���K.F"�wW��S�ȧ�'`�	!�\�`��keM����R��&i��`�'R��^1���w��5ͽ�\l"�Be���3��� ch�ip�����$W2Q��X��H�s�!2
�3�U¬�lX�XF�ҘL����^u�رֶ%b���>�!@���^.��bݜ�οI%}�+���DA�#�i*g�{1�#��Ys�?��|U��u ���)O�Mؿ��Y�����Z�T�M�C)��9���X>����cKV��|��Fp3�-KI���|Q�*4D)f����W�ؼEș��t��-84_�q腟�QdMp`�A׍����`���[,`d���b�30v��%���d-���:[��	`+c���̨��B�zd;6�i_x��c
���쥰]�&�9���v��ti�-m�y��� ~C �'2�������	�� ��LG��nĄ4Լ2K�K��O|�Z�~ȫ����{���/i�e#1���z*���N��l(�s�VZ3X��k��߁���`�7�+��������?��T�u^�6��I6�j)�j�Z?9��B�Bb֋�ѹx��"F�%p�n�w���^�+�V�O�/�kc�Ѻ��+�L�p�Y�T<�rR�&�i]q�]�ִX�h�
 �� na�&�=�k�����^E��P&��?G�7��xJ#��=nV]2�R�9�0
E�)i����V8�`�Ì���=�����0[H>�ְ�4��%:�;��LǑ0�B� m��_om���`W|YS3��^TZ��7�>�3G�J�0��1W�f�{"ʁ����,���\^N�L�fhk��3�U�mO��ʕ� ��)��g�45�D�j�S����j������@�Q����%�1��7��B��ۚU��@|�bϷ�U48E�|(���uBS������l^rEZi��
��c��=��r.���\� �dF�����,I�&�c�6��y$�Y��P��Ų9��#墸9���P�ZJ��|c|��7�	��;���nU��`��O���y�#�wiew�6�%5c�`{X).2��gj�~�J��B���&[O-A�3li�$��:s-����6�����>�� }���%u��Da�l�&��p��WR�d4R!	��~���}[�dUaT��O�5����J��Oxz��P���.v.�z�\�Uk���G�l�j��%]�̏�^s�����F{t��b&+���$Bˬ�"�������Q� b ;�x��*�O�~a�VT�tm��c_{��"�H�	�Wvć��i1�4}��ֵײ���u��F]�l�!�	�OS�
�V�`��!F�Hʤ{���t%b�ܘ�[Ջu�M:|UY	�n�����	�"�?��7�N�~E59��	1&ٝ���u�FȧX�"#1��:���p�U	m��hiu����L�����bvlI:���Z/Z-z6C:���m@vbl%p��貱����lų������Nf���[�M�%Iy����Iu�?�w�(�S	J��� (ʈ��ϬL�����	g�k�?x�ū�h��]Ql���C>	�
����]�o�7��췝��Y�?Ht��Ý�B��(��W�2B'����͙W2�p,�'�'��H�j������ T8��ԩ~��PU�gѹ�bฆz���_���@�-��[�$p�D�a����F[�Jc:՟��;�4�4�+����rC^Z�|	�jN��/{�o@rԕ�r%����DزO�8�U��<��-P@Y"�T�/؃ː.7	�M����!�<�P�5+�����MN���PA՟x���M�v!�)GG)N�К�"�ǆ6����,�wͮ�\P����#���ԡ����M/�8�_��,�[xȁ/0�kռɜ@�MSYR�j�B1>pm�*P�{Ax�U�|���Q����� !'�^F�!��w��)�P/ys�srmc��w_6
&4����1�Q��� v�/��E����.�$/���B�
�~��V�ݔ��DV?�w��φ����3�u�S�����WTL�����䌴���m�>�bc���RX6]J�o��y�ҹ-�Q;_c�iֽ=��%M�vG*����e�zMUz�g��6�X�$���-% � SZKX�E���1�������
�7c,�OpP"�Ԃ��X^Y���*ĉ���4y��^r�W��˥H~�H��e�Y�q��aa���H�Y1���*z,!�ɐ�QZt0�=�_�/�� Ѡ�^w���i}�8��G7����6uuh���Kp�~�Z&�5S��F*����	��>:�/����D0o��AH�ˇ��7.)�G��9 �
�h�j���뾇���Қ�SG^��>3�<ZXv�ǉ���-kFP�Jy��aٛ�P駦(�KH�q}�">��u�;H�V��`���Ԙ�k��uޭQ'�Y
���^�ϒ_��n-*	a ��wۂj�`0H���b譞N#m��%�ˋ�]�)��� I�}��^��v�^����w΅u��S<�w>��3��s�du�ܺ�$��Y�/EX����-���2��V����l?���`��OƺɁ���JOF��2>Vk!�S��ȟL�;/V]��ͮ���~����@D��h����������8 ��C"9o��s� E�uB=����#��B���xe����T���R��|��hV�=b&�O�	Z�5_�G�dwvbv�۴D�]���n�����d��1@�Q���������[��H���&}��5� �{s -D��r��9�B��yt˔��D^b�6Q�a�x�>��4��+H�Y욨�9֐n2����#0�F�U�/��t�N�h&�A#���4u��>����F�2J;/��#n��q��B�=hr�!�f
ʺ�Wk��qO&_���O�8����4��MV�Ø��Z�.@/���j��ۨ8L�Z��[2��-	�������Ke������������F�.�m�=�����G6&��[�HG���Ț2��� ��4�e0L�&ƛ���	�^g�q~�=��<���g�c�f��%���a�F����ć>��U��wK��K���Z�����o���8Oا���4@�)���wv��1�\E��Y����?�z�~�ɍbz�2H��������<�ҁ(��-<0�S�7�@Jh�_��|9&^V�e�T���e`����1�-p��|Ӏ���P�6�����7��=�/�u]�]PCa�P��,�3C�Ne{?J'� +w�Pn�� p)������������54�ŝa�f
~(g����E�����v�Ԧ��N���DN'8�/f�i.G�z��7e��U���}^?��c��\�w��q�g�>�9��WU����I���Gh��
0A:ցR�8n�^�IJ7>�L�3�5��1�n}䞿�����te.�V�:%3���-�0'Z�;A�Ϟ�<<z%�A�4���/��d���| �7�	[%u�v$�Hs�MK7e,�Y���0����ph
P㶀O�`گ�Y �\�l���@�k`��
38�S7T73��#��}�(	������$*��v�QC�M�ji5����1�T�&h������h&/�p�,���\�Ռ@P��Yg�6�������q��-�b�Kr@�˒�E�[���y� �>�'���V14�<���a�cCJ�p�_���ǂ*b4%�6ޘ��V4/���T ��n��J� �$�������d�����޾;JUn@�tƱ<�K-�B��F����F�hNY�1�R_���d�Ț�RoP��p栎����\�0
��1��u>X<��XM·=�����)�q�"�$<��~�<�(����"輻�Q����K��	ː�i$Mq�����	���|�a��ͲK\�!��/&��y�F���n���D/����w����q^0��u�SZ���d�p�4�sa��_nLD<�'��TxMZg�_3{�����!�g;u�J�������75��S܉z��PgZ��p~�:�5o/:��7���5\w_�~�}"��$�k�k�f��rTb�)���C�C��[�/��c͇Rԛn+����q�idXu��n'u��H{�W�홹��$���D�i,�C��U�
��09�殛*;C���s����©�3:-��.����nS3A	�r<��nJ-����0u)���(�e�D��Eq���!7bkw/3g&�]������?�Z�.c��P��
��/��>�&��S/K{�6~�u O; ~�a���0ǁZ:�+�~BH��N�p�Ba�{�A�wV�N>�٫��˷U�	y3��@��qtn#�IĊ~��(�X� ��3\
׉m��?�����������!O�&*ID	��T���\�;�exX@I-����=��/���n��Xs֑l�у����R,v�Z�H<9�a�jwN�6��K�B��	��^/�z���I�T��wA���b���k��b�ӿQ�>4�d��9�#���P�x}��Ai��<�W���fj�`n�@���o��ZmJ��y�����!a��m��i�F����E� z�����kz8}��-�b�Tme{�?=
f'��-������}�E3�F�i?���״Θ	-�����ڊ���*���TmYn��|�B�S�
����4.Fsd(e9mW%^�d�[ͻ1e['�>�ws�l@AI"|�na�ʗ[�m�rP3k,���3�f��S+_�eT���-��Z��|C6i����;���S�_44�/�,1�W���h�]X<��ml,D�+.��,�����į��\0�1&}|�Z���m|@��\9���v�3Yն$9��ǜ����[��6�rx�	܋���X�yN�,bڋ�&�Do�U��)��"�(�㒩xV�@z����r:�"ή	S�;�Pڮa�۝_�J���R��6d�8G���^����e����[94j���v��7m��ÑLy�	J�DY���<fMA��l�-o�q��r�@ �$͆�H�;;
_�;C���Y�6�u�2��/6kH�����!)��2�[�hM^ �X�im��ln���Ƌ�ĸ��~+�|e�r�*�_�50�|SD������-���B+B�h�B�q��w�e4���ŒY�����D�tdJU��m,�I�0�[֥��tD3�(�;��!���,Q�Z��7*yH�
� �S��&�|�x�W���eK5R�V�䨠�!l'�$�h����K�w�}�B������ȋ FG
�3Qp���r���zΏx��Uvx��zT��c�LŐ;J�e��4�"�<�+��&��{�Ի%���|�Hh͉h�  .�,L�<U�{�$N��yi���
>�h�6�r੤I���݉��i���� �k��0�^��-w�!��y�t��ΤM��ft?=�MhY���-,�'�[�΅�&*������-[����cNS��#�2@�h�0x;�(y҈*�p��^n8�I��Yv���v��3�&z�kU�;;�����kX���8z[}F\��&��c,;JL_���.�i��x9c�c0)hI�{qP���"��=���\z�"���v�(�-1X��³h��5��I�Ya,w,��J�&���Wz�h�����ڜ���S�qF�7|fMʦ��SNAl,�����Ά�	�,�9P���r���ظ�d��m�����N��ㆦ��Vcf�n�SE�����R�xsn��.���A1�$��7Tz��#D����ꗳ)��7�?�=yR^�("��U�%>k"x���;~Y�t����a����)�A�w�C#��2�	�[�2����oȅ�P��*eU�� �\��-��0��.�fL׫U���ȅI�������mV�|���J�"�+�����+2��a3c:��o�N��|n��V�4��s���U���͌X������A[�@
8����l�~	�5���*;���U��KT��9o��ڪ���Y,�bF�P��J����6Y<ˮ8�(}���=<.�ǸF�m=��#���܎_46�� ��!�
������m��ab��������& Pǆ�?�ż�����A�yV�|��ܘ�O}�W,>�25���I�3N3�l����
���̙��(���V����pj�\�_���y��t&ꗥ4_S���G�y�v(*����J��]T�դ�_ _�oxe^���� z��F��m���\�L�^���W
T� ���Y����C��:�I@L�5��=�ށ(�a�N�MW��d6h��g?�-�m@�g����<��Z�3Q�rj"�����(��یp�Cp�J��x����pۿL 3�s��i�OB?��wy�%o*�����jw���D������AD�GW;��o�>��xe;�m��d����ռ��/��\�;��`�*��}�����t.��M�`\�j�j+O���rq�Բ ���ɥ�_b�1��9q�j�ٕe�U�����5z9�(������s���Ѓ=M�zc�Cp�E��L_�!����`�X [�����̮���K��1a_=:��UY�P"�5vGw�`����t���D�I�<�|�.�A��Ŝ>�;�Y�e1ʓ�G2�W��� k�Ǹ���C:�4WǍ�0lv�,��P�"��Z<�Rr��B��*�ӮX��L1uբ�r�A��52�h=l;�!�O$�[rm��n��Y��^^�I�j���5r��� A���҂(Ϥt'��5�'8�-���n�)��l)��L��LI����V�ex�ٻ�$�Z�{�ii^�ƃbM�[F5�N�j�ys����>3��5���
��"�P�U������a��������<y�qҮ�ada	 �	�Y\�{�"鞡��E��J�*E~��@<�aC1wZ��@h��9�*Cw��p��
��|�������כ>=/K3}W�������ɇ��(��$*/{�>�d#A3���I����e�a}�Pw7LO�b�)[q��M����#�ă��T�l�ԝ��߸Þ���q����&�� ɇ]���	�Dx߭h|����I�/�72���"��;����_����].C(�gn>ȯ����w|8>���H�,�\`݃�6T����m ��	d���� գ��u�o;��}�2l��p�Ę@%��1X�lk��3G1�i�I��W;\�\D�����'���s��:u~R�1�e������O�hlF���z�+͹����1�M���!2y\>Q�d���q �F��b�y��꺺!5�TKv���Cu~�I `�2�����{�6�g-z ���Gd�2(��P۽��خ'\7�4�̓`Q2TXӄ�B��#���㠮������X�ތS��0�6a9JZ�yHU(/�?�Nn�LAfp	 �>���w8�s��$��	M�ID��1͚P�Q�����hC*�fR��t���=�ux�
�j�V~�xa�z�L�;��yV���3������M�Xoj� �.?k��P�YT���vYPqsW���;�Ly�~��pxLܜ�̇�$ԡthb0t���(�4TC&�|�U�Xz����3�N��\w�^�
#r~��f�|���L�П/]��B1(���>�j��-G>,<��!�r!��]��l-�|wۙ��1�f���~�^����c�^t#Uo<��R+0dD`)����xbX�l +5X5�E�y��w{�"�i���K'*�� ����%��^2ɩ;��)�P�A�"�c��LK�lc��«�
�G�%<%���+�R�o�yz�'���,�_{'�?�\��\�/�ۼ�J?6���v�i���I�J��c��S�7�Ԧ��\���a$ܗh�/N	�+<�n�r����@;t��lʥ݃��Q�bbWNCvR�mV�!ɘ�����L�f�i��/b܆�����7wr6�h6�mޮ*h���'�о�za��s�.��B�X��h-�|%T��"]�����((N��*�֚��=?$��q�S��/��HE+2+bz�s�8yd�7-ed�~8aְ֒�c�w���3N�\���c)��KA~�o��� �m�F��o���CWB%�=���I7㮒W� ��3lUs"������I�/�����Ҵ\���m�������)�J*�����@��1�e<��Z�bt&�,l����Ig�ڔ�7�( �a��$哊����d�mqu�00v5ɕZ���&n���/4h.��hC�|�C�N�7�{�|b�����L��ޟ�*."��#��fף�J�55���i�ap�G+�zĕ*�
���<����UQ��e`��SA)ם�$�(�/��H���4�ʔ:�IC��y���p����m_��H̊N��*�<���H��-�b3F�c�
�PR���֠3zP
�q��Z�~��N}Ѳ;���qi���ؤ�XŒ��g8p"u�O63��#鍋�oo�R�%�E�%=a����EBv�"�H��Bk��Mg�vG�h�1�Bt<H�-}h_Qtե���2�mh:7�v�G���~��q�����5?`H��o(��H��ï����  )$a�4'��Q�!`Y�t��<�GL�K!9�q[ըU�8O�DVd�e�@_tǡ�ѐ@����Nt4/f�-�C��w�q����i���Qm UD�i�������:��#����%Q���*z[�#j^-5
��Gp�#�c{Ej)ju��2�15378IAq�������:��Y9J�g+�8�$��߁��6�f5��KC$	�������i��� uQQ2�_ ���'s�X覡��'ac��CxV�����JX�ͮ�}�C����:���5��c�!A.%ӿA���U1�iH �R��Ի�3W3P`T����i���Q���Tօ�6��y問���٬���h�H��6�FH�Ŋf���x���o��5}&W�ǃ�d	��g���J��a}O�Zg@�� (�pbX��+ R��f�t�}%R�)?�l�f4���3�)G�\\.Y&�F�� V2�%XR� o���i�CZ߲���h��HWAKj�bB���Q���3I_N���.�<늽c�Q���r�}�
��l��i��e<���qvm�|��>M����F\��I�<�0v��+Y=A�oM�v
�U�<u.������OH��Y��%�ё����^�1<^p��w�H���U.��7�¹gd<��Jx����w����'�^F��ԧP��6�Ǳk]\��y�a��C�oЮ{Z_�>;i������7�Ӹ�s���pu.��-��2�T/�8"��>)�I���(����/����t��x<�$�7�ݚ�R�=��}�}�����'�?ǹ~17pY��O��T��`�5b��04��G�3z��ٶK���#�K�u���-��YH�7�T�&�C�������Um�K� ׂ~�i�n�$����#��5��yO;9Ԇ0�P-�.æ���gQX\.�}�����l	��ltYO�k^�	��p�P�dB�;���jo���ru��N�bǋ�Ǹ��ܸ�7�j��x���9���E���#����?�I�@Ǧ���L�P�hmo��7�<���.�0����oJm���m�ͪ�}���ߡ�lP/�,���y�P5���Or�@	TkZ4
�/eE$�๦m9V�L{�8�-��fԘM��Q����]Q�2���������.|�r�[{�ۿ�~���<y	\\��E?�z�a���̲�Vs����R�����P�cC����eW3����(�Jwv8m\�}u��t(�ѳ����v�<��?��ǨfÁ�fis�2b֚o�����-A���g���I���#��\����s��m_2��pv�/�ڸN�(��{�2�ŕ��<�O.�V��,p�-�J�;��N!
:ń����}���������������̢�"eQ�XRsն,�4��ӹc�Wl���N��2��̨���t�j:/jډ+/�q�-9�Є�������E����$���r\AEs�R�V�lߞ~�1#c���5�+�A��Hj>iE�׍`;o� �pܯܠa�@��P|�K
�|oP�2���
z�`��/��VI	�riPM���m�oWZm/
~K��f]�/1��g�����_���������le)9�Eۄ�`^E�6i_��N,	Wǀ�݉`N�D��N��U�(�́s�-���V����t�A��I{>�؞��?ҿ�0<��3爄�Kwş�ȏ��>E�|�R���2m�z$��G�6Y�M�v��Q]l������k5�6�.�
��=R�D2�C�� �vǽD��{.G��8�ľ��l_3,n�f�>�*;���\����5�����L\O�@�M=kE:Xs�<���]�7�;�Y�����j~�[�'9ey�('�6XJ_����&��,�;���Q ��~m��DI�BZ���쥐x���ʑ�d�������	/H?�ٛ��/�m���;U�"�	��ł|>=�I���åh�]3��1*{���bgߗ��F�j_@���{���8D��]o�l�_fI����w8@�u=���@�'Q��VWi��!s y1?E�*����\�i���?"�J�l4�U[,J-�A��s��9��ؓT;m���/�4Q��G71`Zk�F����O��Ӳ�Kk�h��f$L 	������8�0��(���<��Ѿ���+�1z3|�P'��\�Q�_����+a�ő��E�VnG$#[�\�z���U�	�1řs��dE�n�L����&0P_��u �p�u;&�P[G���@KY���6n���uV�r�-���#
�X6l�G��W!��8�q���YT�&*1�i�����vlP�A)֛�qv�4U�T��A�rʍȵ}����S�c��M�B��\����z�-S؏�|�i����Ug,m�u�-YFz�56�&Y�U痤oy��Ź�Y����a��� �=Ѓ��+��5bi��ش�-`X�o��.��߁�{��6G�U�������iS����K�|�w���րu��maypؓK0DU��j��ta��]=f�6���e�Y%�?��wa�Fy �A���Y�g���^��(���EY����!�ј=��'����Þ˯�Z�"Bo�Dݺ���f�x�	q���4���yail�����"��p;�Q�r����%L���_�1�����G��P�0D2�V�h��or7�=��bW�K��
��2�"/*�"��0���
�G���s Z��!�c�4�Z ����;I)����tqwi��¥�Ѿ+�j�jy�R؞]~�~J���7_�L����U7�,��֣m5m'Ϻ�$4�H���~��\}n:�����ϯ��Wdt��<�{��'y���01CK&����e~�"��y��{��͗�|μ������-��&O��,�qc�l9�&�ND���ɽ��kh���%-ces?^��SK���9���	H�K���3��	�G���v*O��Ɇ�t[���wh�a�j���j]���zY�}����2��,BL�G��&�t�u��D��0$~��8��R'�3f&9�k�D�h�!㨴�;���>�B��7��Q��?"el}'㟿c���jX�h��0�>J�J��XQ/Y$%A}���(%0��,<<:J!�!}���	����)~�E��� �����Ŝ��诚����vO�K�zA�#�0$?��Y�!����
��|�`ϿV��bv�!�:Rm�X�1�ø1�v�����@x��}�PŠ̛�Q#�����P�1��+�Q|G�1+�r.�i]=�&�8WdI&t����ֈbDw�3$�R�#�='��@e��Ⱦ����<���L(��uuV"!�[��«���]K�����f��`WZf�NҀ+�_���[m�?n�p�l=3��u��Ν=�|�\�H�|q���,�`��f/C⃥/��hÈ���Iҡ�h��rW�US��%���ӮaN$��Ѻ�Sn�L���ӥQ����](�.�a\Y�(J�� Nx[{.��g/!����0��2"6�3��={��)˃� #�9.�b���P���8�Y��f	mF4�G,)8�� rӊ�rI�N��5�j�m� �^Ҍ����wRF��aQ���tC.�X�Ǖli����D���|�[�f4��D�ݶb'�7f��S��1�]+�{r�����
^���OI;5[T2t:�2�hk����o%G(�O*��x��G�?[����,�*(-9%vx��T8�_������:h�E�2�Izh��I���fw�����󇃡��;�'�O�/�Pj��}9���:���&��G�8� 1fQ53�Oc�#G��j}�l����ڡ�ѮGd����G��2/W�+� :=�L�����mq��W���JV���ݭoeEء!B۩�X�_�0�����4���WaY��1��=M(J7����`���C+:M� ��3�Y@�ap��4����&|{�Wb*�e�>�]�s=5y���{�G� 9����@��,�/��/��sd¼�h��Ԣ����I� )]=��2�.����c��sɠ�D��T��.�KJƎ%~��`!���YdQ̂�&F�r��)����>
���1�O� ��;0���~�zf){����-Yԙo��D��5�# Y��5Kҿjs�F
T�b�ho/���ҙ� �Ķ�hc�v����)��;��`�'���σ�]�u�O���E�^�s,�	�R���{�T�m�A����MK��������uZ�jf�t�E$=��Q��][���P�Q&.x?c���!��o�c�_
i9%�`GDL���r�mX(��%��:f��P�����r�9�>��U���k�><Y2�*ƈ#%�41��}��^��uR�R���Y\��1EP�'7�����.�d]<��m���%2��jcw�������9@����T��S��{ʊ1�na����aj$�m�"3�5pB�.@��b���sJ�l������������@�(
K���t�U��_ƻ��i��B��|��z1~�>$טc�.7l�a$Z���k�4ڿN#ӝ���������R*1����	SDQ$�(�5���^u�_'�{q�幋�K2D��ʜL�/m�v�u��,�����Vϐc���sG��@�f���H�o:g��[4n�Y���,��Ƚ\���f܍�8�=<)}�,0 ���{9��(wYq�j��B���L[���N����/Lk����Q�e���ӱf�#ԾKyS�]�Ф�w�{xH1|�}IA.`�*|@�Qjz81��Dvs�Iħ�"�Z�g��V��+����CK�D̅ �(M,�R�C��
�W�0��y�Bl_�a%a�Iœ� ZG�UX߀���Z Mj͊��=����`j�R�4�����g�n֩-w\`>5EK��,��װe��7"y��2��:��S������`֙G�����Q�6d��U+��Y�-φ�:2�"e���
�GC��B;dይ}z�A�j#�^��)f�f�7�
�8��/O�n���u'W�=͖�)3�RD}c�}��0W,�)IS�;�P�'���0{��,� \�[�:�A&���ʯW?'�̎NJ�hcS5,f��+O���(��[ֵ��\��XU�	@ݶ�c���y���	����{��r����x�ï�p!45B}E`EWr�E����0�*E��ĳ���>(Mag�s}!�
�u���ȳSq�~�-h>e��%�ʆFCg����w��̠�b|�T�t��~�Y*�
�7�9�?:8�S�8"@�:2՟pI�%�/2�	�[W�pL��� �Բ���6v��E�C70��op�I���
}��_=�sMCqF���]�B�}��!���~���TH4��$*�K2�ڐ�]�΍Orf���a��'�FDr��	[8b�8�ad��k���Dߨfq��{�B�VTt|VL��x��V�$[F�� �YD)3A�pZ ���Z�pJ�#��.����+Ȑ�����[�U�%����a{���D����/���q��:�TB�����R���eh� �3!�f���mvs�eA4H�&��&}��OaS§�D�N�I�r���0�j��ଁKF�Ő�k��Z.����W%�zϻ,�>����]�O'!&��3QԴ�RC� ۻ����=B\�+\G-���s��P~T.�)�� ������_:��KD��'�0=�ߜv6�(����g��>�' Dz��K�nY�6�.yM@Ѭ�C��+?*��ܪ�(4z���u���t�	�paKcUNyW����E�&�Q�O�S�h,HĚ6
4��C����OJ�)���w-&T�HC�`&��-Dv)���8�+U��	��d�k�pI4�y��Q!�@�(⪼*���r.f���.�i�5�!>Op��r��۱/^'�=g1sd���4��T_ ��M�MU��6E �2�򈷻Q�O�֓�b<g>�f:V^�ծ p^��<B�m}�c�Cq��C�-Kd�)�d>�6���/┳vο��=��)��4Yx�� ��E�?L1D5��G�R�QyEr��z�Ǯ��í�4��W�����q5�I�PR���՚E<�iLK�f��Ȃ�jTGZ:m5��J昅5����K�{̹��Z��������3��_꫚�/<��}�]r0Ǹ��i�$:�3��
���{������f��M떘u��m��"��J��V�`وG�D6�07f��״OР�Gf\��(8ؾ1�%�s�N���h�b$]�!���QX��k�(��
�.0���Z
l�����tOj��d�wց�g,Zd�7�+�ӈ$���F\����}�R�����|p9�{I5��W�ib�����S'�� �H�S-"z�d�~M.�8D���4*�5�v%k�Q�ջ�h	O!�Nl&dN�����\Y\�������i$ ҟ��=z*��ϖ���Ă�iz��ggl;O��L�A�{z)�g�RFx�	�D.�3VAp���cY�󭉙PlZ��`Ud��G��)�H(��+��J��:������Pw�ǒM����FxFI�<�{Q��)��M��"����@*���"k,�����%Um�����02صS��t�%oWb	2���j��p�Զ�'%4چ���+�ʸYq���z��� ���l�j�8f,�D��(�?~~�~<�7�x�Pz��0o;HZP�����������E��L�C�� �/��_ѧ��2k��^�lOn�Tq^u/�bZ����'B�0�|�	<�mE�V��!ϫ���LV8	���_��	�D�����kL]�,��8Tж��2�ԗ��켤��v�+�]Kc�i(���5<|GV����-���?/*i ��e R�����I��{����XN!������NA�Ьk�*-��<qI�@������G��	��W��V��"���f`�[�.���P�9�p����<~Nn��y��,����X���4bUTf�����$u�O@�/0�Q��g��~}e}�i����٪g�}�cUZ��m�E'�G���`�/i�e����Q@��|�vw�S�����ĉ	�ח�m�C���]H�?��6M?�9�c����P����R�8 ��?
cR]���<��9A[�*qL��I��  }�lW�+ƍP�k�{����[ك��'�f/�X}oUX��
X٥�$��8��tj.������#b٣x']��y݌�:ZU��W2�%C��n�fև�ڗfm!fE��)e����j9��d�V7i���� s��7Wz<&��e���4)�_I�I�R?�6�)���H��ic7�@y[Ϙ�'3j��
��Y�]�"z��R���SKe�d,�����V��
5Uj4���2�F*|x�w�F�H錁�8�MA=�E��8_�y���	OZ�˹�b��2��x;��b�oe]��u���p�s��6��b,�������Z��
�3u��n?��F -R��?��+�沲p=8�oHaC1!6��R&&H�����2SWt�aH�=+bE��a"���icY
�������ޤœ `��(��|D!�T�r�X4Mwp�>k����,�Z��6qۙRqs���uM���<�����?h�iUJȩ��?f؆�M.�=�Z�h^ə��Ec߽P0}��J� Ot�.]�
����hU �һ�*�~�im�yO�nŲ��~|X�@7?�����jÒ:h��cq�(���p�������%�m��xbZ�����TB@�f��1�C[��+ٺ��r�C�K8�9t_�^xl
	��X-&�3�p�hJ�  ���8l�����F� �-��SVH�1�t	�
|F/���{"g.Ccú��{}�� ��U[��]E��B�Hu�����;Q (�̆�Xb�`�*�W��8Ua�IBT�L�&]a�]���+\�{�ܜ �Ս)���~WLQ�V
L9��\Μڍ��1�"��+І%Zs_v
���5u� 7�.�9���I=��Fњ����c� ��,��u�\f���-�m������*�W7Ǻ� ��v0&��R}.�X����'��(��z �52� ��dO�G����,f��Ŀa�(%A��pƔ/���^}����Ua�q�j7!{u�*�ED�A�߀X�߲l����v_t��3UߋOWN#�s)�V% ��K]c`��Sԁ�q��\�����3h��T��%����.A���è����?�"����V_���M�쾖=-���gZ����!P���]^�m���P�d�Y	�k� 䣇- {W��7̣]����_��4�"�d�����T�O���uE����=NȚ��iK��P�aބx�b��HqK8�7�h4a��gk��0��2bO۶q�Aùp��1j���Y�k��r�,#�<'����z\.h����8wm��ܰ�~
��Os�������}��o�����P�#v8�&$��7K��*��[��#bnKf�U���F~ ��h� D�M����D�QF6�`u��}֖Nx_3~��xb��jI ��{�RU6��թ�0(���6�Bn�^q����}K��}�^�8ZU&�֔�@�{Z��t����*�o* �P܈���o2u���LQN��p$4- 3����`�ے�����LB�(��!J�!k��p�>-OoK�I2�cy�����a'w�����|G>���]��IK
��4z���(��6��!�b\����$�ҌM�L�'�y�B-����0��=�22��J��:H��c��"a[/�0z.Hp?�~�%�!pȑ�qGP6+�d�b9�� �� LK�LwP�gr�^�=�I�*�Һ.���%����+h��0H��H-���:�g?���Å/���97ȕ��nqG��?��:z��
�����kj�%[`�㈵^�f�P����]��P�H]���t��5��wȊ*B���-��STt���O��������`S֢W=�����d�u�I]�L#mt���d,������!�=OP��kUhh���3��� -�(������6X�Ů3w��(�W�YpV��J��Q��%�Q&-�Q6�u�E���K)|�u�2V�[9�Cϟ��wE9٫���%:ͷ�.��]�\F��S>��튶Y�'�_خ����e���d�@�����gT���%��
��w���y��e�ŪC!�Q%��r+�V�s�Գ���� �YD���p��,�,l+M4��b验9B�����-)�A��7u1]e$v���{��`Q����%q�RDo��ާ�k+W�'���(6Y�D��Aָ�e�.��T�5�z@�p����^� ,+-sr�Ȏ�g�l��rOL����;g惇]K�̂!�Ϝvu@����j:�u�졔�"���p��������^���gt��[��Y<�I�9w،͜�X�0����0�B�Ջ���"�tȑ?�K針 ���Ѳ�H*&NP5��^��Al�HH��ȹ��'I��TL�ʉ�n��?�W�����u�d͞�g�k�| X/"RGV,y.��upgؓ7:��{A�
��㕜�-xt��+ዋ�rס$�,S�����h�d�s�ʸ�"�;9��v��J�t���ץM:y�X����ܭ☿�इ��6�{�b���	)�u&�|�P�-&�@�j�\�:�]g�]�dWҍ#��HQw�����ф� �h���C��38�Ӥsiٍ�I�/��ϵ����	�����]��>�͕u���-,e�#] �z��b^����SI�z���|/��M�=9�qX����L��'p봶mVM��iϞ�K?���,BچI���xd���6��ގ�c^��ݴ �N9�c�!$�4G�)MϵjNEJ�$�a��H�NA���W|5���%o�B�׎�$���\w!`!�:y�}����=t5�y������-�;N�>h�ʹR��n6ѧ���v��;t�,H�!+[K�~XZD���L&DX�B���'X��A D���P����r7�r�]ME�hO)�[�}�x���I'�$�i(�v`��Ld��7 T��E)����xC`F5�x��g$���Vy}Q��o�|�i����� P_��5񀧽���z�=,�AOp-"�������kE��m�[�Y4�d��;�E|I�eD����(fv��Ƌ�Ir(	%�����dARFl_:*i����H���ngG��WU$�hZ#����,�v-č�*�{,�)U�������%#��� ����ME��dH�eK���F@��j��.���.��6����Jk(���-f`�_���@Rˮ�T�/W~�&��E��69q��Y��?�s���r��Q6	ؔ���F�U�q��W�v��{�F*�A��n�vU>���\;���#Lv��3���
��WoU��!���[�q��R����=
{B����V�ʼ4�lx��@���U���X����x�, �Mg#�p��N���n,�B�����ƕ��	k
�1�5�D��K`�5���&O�_�}�W_t�#�~.���j�X�������i6��^��mL�yu�o�8T�$�E��l��'��	�)�Ļ��~ԛn%Ɣ�R;�*� 1�LX;NZtym߶������ ���3����y��"�Fi��`�z^T�S�z��cVn/}�'Ip�+!��y{Q��&�.�b"Bu�9SI>���/�Bڷ I[�('�eH�(���)H��b��	���+�P�w�K�$|��ww���F�]m&X��,ŝ����^q��Ub�I8ilPh�&݈�g7��"-�W/���ҋ�"�����J�l_vs>]�5�������x�O�D¤Cj847��e�8�m$S�R�H4Ř�o�' ��I������)��ӾP7=j���DX��4�z9�Ņ�����Nu5�$n�Wu�4�]�C��h��J���|R����@�n�*e�EV���j�Q�!�}(%<������آ���$ݞDJ��p�h�Z�R�r>���ݥA�:�]�h��C��=]�-M�]���(4������6�F�%/���`4��ԊA	���������ٚ�m]�*�f�3��#���5J����/��ɟ�d���L���.C�-�W��)��ʥ�\��uh�=f������?�V6/Ƒ���e��[_�l�m�|�[�cذ���K�Q�_D�
8�� Ⱥ^�U�KK�9<����;�>����:���?���}�Aן��=�4��F6�Y�k9���i�H�)�&��e%��AVs�x�Md����U���P��t=�6��E��N:qǪ�ud���QQ��$?}��l�Xs)I)rq$}W�H�����*�����6���:]��ٞ����F/P���Ϛ�ܠd�Ɋ��U��j��vO@ɴ���I8tw+�r��+.���	;�7���cQ.�"�E":��w���1�!�v��Hs��ZHdL��x4(��!Jfd_&��ٱ̌�i�1�K�S'�b��-�Q�`��s�tHW�'�`��Qt4�01�_Rݓ.�L��9�ɑY�|���⚫��q5P��v	A�U�g���Y��h�`	�ᯣ-чl.�GhhU���<�_�f�����+됇ن����W@� ^�2�*��jG����j���Wv�.�9����hO��n��A}˃�Dd����3/@3z�\�]W9B�$U<�U������ȑ��᭜�����@˭Z�F�<�e{���2�(�5�C"'[��U��F?��#�PM����]�&����<8��wbLzAŪ0��5�f㑗�hڈ��.�����_*��+P'��|1�`��LO}3T��:�ZP�,�j�h~7��f|��∪���_uΫd��ﶘG���:����wˣ��,.��Ñ�0 �$q�\)���nہ3��X���9�˸}�?�`�E���4_4h5�`�V�!My/�P��k���y��!Y���h6݉�=�_�_0bݿ`�}=��P�:�Ap����Z���
��S\�E`C���*�P,��?�P �,���.��v��>Tk��e�9λ�uu*�G5v�����<����Ey�du��,��<1_ۅU�'�Ii�]��(��m��;�;���Ѓ^�*Z7GeJ����=��д3%?n�-m�{a�b�շs#�Ʀ�6kR����߷j���ZuZgj�&̻)4�`���ф�X:Ao'�[��F���὾lw��qj��6�d�#�������	���*�U˾F����Ew�����i��o���Ы̿@09�ۈM�b�$z��>�*�E��C��\��q�&�1�o�SvV¢m�/B`��naF��,��;}TL�����¡kkN+OGw.p�s"n�n�W8�l�[��w�x�b� C�>�nB|����� �+�����O=)6��
��'���m�~6�t>
�WF�21�rmɞ���;���Dd"�tI�k&�����3����^�[���-K"�f���� ڎ��|�ݐ��b���/2Xe�E,5U���87���qfHT����Or�������'4�;�O .��)e�}�^��r}߮���0�HA���L�dB����m�TVZ������J�1�ݭ��ؤG�\F�|�c�P]OߺrV�R���hf����%N��������q��+_���;�#½��wQA��k�Z3�Wx!z��N`�J�|�ܸM-�U�y���l�Dޏ?A>�g�ԡ+�v�˫)]ȍ)y���yOl��7���O[��V�1�"E�3���kZ4Wm�U����ђ�(��"�����g!,�Y�
��[�$Z�o���D������=7��Z��gɃR6�H�!�5Z�t�������wT�`/6ؚ�,�������I���XR��^�����cV�"j�1�Zyv�c=e��a�N�/1��U�ն���Y�\�vcz�*�i#�E�9�1��55Y�xz�6�P��z˅Qg�2��_:�$P���U���*F�����"�>N��?���̄a��1�M.�p���٠���o'�K�rN�`�ʋm=�I���>M`�_zy&@�=��Q�� ��#Ÿs�p6��+C�7���>��M���+���x�a�)�m��f�`�K�"�G�y��n�����<�*H�=�XK��-XX,h�Ͷ�
_�8O�a=��P�O�ɮٸ;�2���a}��`�)���LVSe-=V*k���[X�r�	>����- �uK$��Nt�n�C����5����f!��	ʢ�`���/ ۞�~���d�i��0ܝ�'E�Ȉ5/.@�S>7ʈ�`�&���q�*}6�� n�}5i(8�ҧj$F;���3�ui�#l�{�e%t��/��;���V��@U��ZK��4]�{ ��+�!�*�1�m��/f�o��Z�
n��f繄�0��~A�\��=B��<�<��V��2&?�̢�݋�=F���Qu�����χ�aj�Ü��iQ�D�X��h�Ba-�`M�Zl��F�)p]\�*�rt}d?�#�'��/͋a���/�������Cj2��m�D�VM��+־�r;�Ux�͟�˦�р�n�t'' ^��Й"�RTB������h��Xci���:^ �A/J������(bwV��.�]�فE���_��-��Es-A�ٳ��҃�(�2A�
�HZj;��"�㮀�w������>��~�Ԭ��o�cs�4F؅��+q���]�W�EQ�x���:�:���3'��ۚ=��@%{OH����H�=��F1�|��k{�0�>�nq�߂�B� �!�&�Ռ�)S��k�|�GQ�,�~
�J��5S���*K��3��a����$�T�r��  ��	��� �\z,��x��^7� R��:}cN��P6��2����z��o�Jׅ��^mS�E()�i�#�#��Z>U��2��9$n��tyܒ5��ے���om��:��&ZZÉ�����g���D�(\48�����{���dR�w�� � \�ē9�R"f���d��'�g?vl|�
�wnSJ`��3\��f
��[���nyG����}��vG1�ȫԙ$�t*���f7d�ҥ,}U����XyH�a�y��}�]�xG�tY��.<e��+F,J��|�J��O�;p�G����%��3��|:iF ���q�W�4���!�;,�Z��	��s��vèVBtkE���I6R%��Rb�Ԉ2\�w�D<�Z����J����-r&���s46?g��-/qt�DS����v�>�6v,"A83��b�o��핫��L�����_��&�"t������"xY�X|o����|)�7�A�ܨ�z��y�ڋ��c����Qv���4Zݦ��%��]�sr��k]�hf�cZt=��l�=\g`��0�b��qUVhۀ��{��g��
��GU-�q��%#%�F��Z�įv)�>��@��k�5���*�8Ow��4�q����؅������!䙠�n]ԅw%frTH���Μ�&pN�PH�0�������e>�>-U&�D�8vq_���8�Q�Z���9D!�����z���8��/�l�	����F�g��;8Ǔ����x����s0նv^"
0<g�99|�_\�O�\��]*����w�ߣ'Y�k;���
���P�ܷta}�C+\G���]�،�k�$��=�H!�-yR`�v]k'-j���/�;IB,�+�^��'�T`Y��q~���dC�wW��*ǆ]���B0
�m5 ץ���iB�N©�@J�@8��ǩ@ ����t�������٠=��Qב�I������Jd�)ͩ,HO��)va����^��� �~C������DXm<�|�SAg�C�M4+�;�8��bvb�j�az�6�iQ�Q�/��w*!����h����mL�
'���e(%L\�"i/��.}��:�)��!�|1����ռ�8Gg����s���H�P���:�e��l�D�3�i�����1����}��#7��U:eӖD�o���{FYQ�a;M�!d�g�EW��s�b{ƦK�V��$gC?�A������`���~����n�h��o����IpD����]i�Α%�nRX8Q]A2�	��}T������a�^%I����[Z.C4&�#�=��~�S���M�T��W�:�%5���0�f�����k\�C���eu�����ȕY����V�Q�i��]=�$�;���l�bXz��6ff����C @ЇP���nO��;�'쌬}U�Wp����#�?N$j^6CX���QA��8�p��������*�?H���CF�"��wA�T����EׂT�
��^�����o���.���������{i� [?-V��+3b,�*��-�^I���v��aq�����mzm�1!�ҽ|͕�J�1�&�K�R�%9�ߙ5F�7%�a�{���cɖYнfLwf�	"w�����#� .���֞R�	h����L�4����&�yG���bsˎ����+���`fgX�O�z�.e���E��`<3��Dq�z�,�bQ�s�%�bo��^��!㩥�/U���cԫ����kQ�l�^įpcp�n�@�1o˛I�*}�Ç��6��(�<��q("�L��XO��/�\ɗw��������r�u�_���w�8�h��� ������Z�k�����y����^�;Ru���� u(�QJ����7WE))����WI���ݴqN�2�(n89P��Ǌ`}�9ʝ�>� #e���P�J&�y����L �g��⇌�b���[)�~V��%�נ�����r��f#351�`f�aUbJ8#V��� Iym�����-���+m1�X{ww��6�p�w�it��껌@�y&�w�S�ҕ���Go��	������-iFnK/��t ]�d%�S'��>�����n�T�c�	��_��Y���j9�mk!�^�t{X��v��� ![�-:�=��Y�#����Z[?�(��l[J�l�ο5v�(s��c���vt�hη7A��z%���J�H�����ܣ��R@�nKuB5��ǝ�F��R����\��:�R,��A]Ié��7�l��>� ���t�W�u(�a��YpC��������d�D�%�`�D�Bv�K@� ������c�|`��4K�3j�G�����Z��b�tߣ����
��)Α�3�+�v��m��cA�� f�W�~@�+��'���	�C펴�Q����)� �.^Ϛ�L�wI�y���ȣ��}�HF��O���@��r����|T˙|0���_�P?z���$x85Q��2D�ytSĔ�_(�?���^���S��>dS�<�!C
��w�)����wo����}����j��}��A���c��F�d뇒�'"fy�tE�AM5�ty:N�iׂ����KK�=��G$��^�Wһr}�jR��X���p��(�%urD����9ԅ:������G�ܩ���}lb�̆F��+VS��H;��������G,t	�~�rʁu6l3��}�沷c�ڼ���:.h�2�~�~`��L�0WK�����;"�E�{���+��K�GK���E��]H��>`~Q`��dB'ox�hb��L�Қ�3a�Kx_.��;S�I�Y��\��F�����y����S�4���RR'-�(�L�r��xf7�ls�������a�m�@`~&s��a�k��;���"�����L*c�����O�nS#Cy"11��i���J��� zr8Ľ�ζ���Z�"Q̛�,J*��!��5�K�����e�ɴ��8Rj3���Ϗw�+>�ۤu�V��c��h��t��A��&�Qyl�Ȑ�Q6����֡�1��Tۮ
���	��X��km�vZ��>�?�sL�xe5�SH�i���ho-{�����ߋ���X�Gu���Ȭ�Aǚ��ń�M���L!�,��H6�zhӞ �ΠI�����l�"��:�d��FH'>B=w}�W���u2�Q����������:�(�@�6{՘d��=U���G��E%���7u>щ��<�w�hcC윈M����TTi{����|x��y,�ƿ:�_��ߜ��s���eO�ꕼE�O���8�#�0*T�[�9�M�K�W[�a�cwQ(:q���c���ѯ�a],�+��-Q�/�g#�:����&�`�uK�`�C��Q5ht�W��bU�x=��Z�k{���mo#�ޤR�N^�����	,�@i���Ht󑢃���ͽ��[�k�5%[�	�u�q��.�3B.R8��=��zg��K�����p��k����F�=��"݁��\�ŋ�,{P�sQ(Ւ��y��S	ŵ�����`≔�=��*R�(Q�7^ܴٴ3���3}�F7��m.�d%j_ȧ�^���)V%��)�ǅ��~��k�	φ?��nlܼ}����[���=��	b8Y��_۴�d�<\`�4`s�~)���*%��o��k����l��0��n.*L�;*�ȥ:P��S���v�`q�p�['�KIQn��)�,�d�UV�npӽ�������c�!b�'�@��f�����#q����D�H���C��ǃt(���Yp�&X�{��׼�4蕬>�]���̢�����q]���c��y9��:�������uog @���l��������0�Y��j:F,N��{�Z��L6oi��.�Q/�qFJ5H�[�CZ�S�G��]�9�܊��[�	�Վ�KK{�1�X������>l��Ni��G1G�}`e:�*�[��`����jy�"v���X�pV��P���)���������� D��RFy��h��6r�\kT�����ʘ���S'�����䌄h�s�0E(�u�q(3'9�f�&W\M*�����jp�v���c���c�d�Q�-K�Ŏ��{/sL�ۥ$�V��e���T`^9zN�.������w�@����⏫��#��C E��-�AمB7ߕH��Ԁ�"V���r�\�K�7�K��:j���O/���J�����"�~k��޿�$�B�_�(�{0�gۅ���d[!��Fc����2 �ߑ,��m]?L>J7Fv�ȃ����Xݷ�:tz���.h%>"��d�d<���L��0���r_�n�\M�Hl�%�D�{w�6�
1���6zC��/���^0��M��n����t%�T�XA��?3���k(��G���:ؤbP,�#���Z0KsϹA�D�Ǐ��]]"y�/@To�[;Sf��{KxF���a$�^:�ߜ-�ٷ ��6|�tZz?�%y�ۋn'�%���{/qW'�P��9�֒	�o���p��XR1�`�:y5�$abQ+ϫ������l��ds��8&��\�x"��0/'n��:��%��d��������(�S�H�嫵���`��!�5}��]�7�C{�Z1����n���d)k�CLp	�f�C3E��Y�lJ��}>��+;�(���_�UwB��x�<����yi3 Q��VU�#��uJ�:M9�K�c	�lwT�z�`b�T59X0G#S�y��W;���O>^��|J *���	>e܅|�f�Q�z�/&$dQX��Ӄ�'9��,�*��%�0��j�22���=��z��6�Fڱ��(3@�Za�c�m�d�+�pa*-s�;4�2-�����S���v^�����L �W�ɝ4�$�
�r�
�ca����fŻ���E]�E�j`[^�1�	8M�DusR���~\�W<�A���f��m3:�qM�N�o�?\K �B"G���ڕ9�S�\���}ҕ�Ri7pB=Q&˾I���m�:���Á��0̹uO�a�|��<��t�� _�o��4�`Kp}kq�wƱ���@�I֚�ЏN,_�����e�%�r��?לF�.�2�����/y�r�u�1��z�_э{:��}ߌJ�3��r�O�{����\}�Æ��F��<iד%�a����s����j��}��ˑO����>e|�>5��M�Mh#��Y��B�H��mn�)S��h��D��Rn��[�|1
 �*�vi�Q���x/�L� ��na5áΊ*�c�_y�<O��Y�-�d�����)���L$Q��1��<���g���|����s�O��ݮ-1d a0N�jbm*t��M��u��~��@�1
"��� p��|���� ��㰼�v�V���B��2��
t�H��s(՞�E�qT8z�}� B��	�,�8q5I�7�N��H;Kd.���ܜ���E�(���\,��aiO��Yp��!E���������(4sc���R�%S���Knzj���3��/<7���Z�e�[mc�<@,'T>��۩8���*1�(�(&�=<�R�������z�mG���n�d�¤�E�ܯ�`]˥F6{7u"Z�gr'�9�A��t,����tI�G!����]����jY���>�����3�DF����|�X���9*��T����H"�PiS�i^�=K-�TI�u�a�}N�jY��Fh����V�,��+�Fz�Q2.5�zH���*���e���
�v�'[�3[��9���Sl.�oy�j�|�ޏ WI���N��^3�eV��^bʿ��s���
 �N�N��es���6u>l� ���;����������?�Fwsc�����}�Ψ�x�˽�f[	�8��w��P�q����]��/ĉ&��0P(�E%�R6J��1�:��;4��K㖊`�B�5YD����o�����e���Ē���(����bW�+t%H*bA��K_\�� �� vp#a�`<�� ���`J�D�Aw����S��Q@ϐ��(���	n���Q]*�[��7�^,�>C�*�1�4�( �zi�I$�L�?�Cj�	���������
*&D�,� U`/T� �.�D�|�,m�k_ X�YY9ZHH�9ц�e~:h&��+��XR����Z���2n������uS��m��ל�ы�΃
n��{����?n��ՙ�YK)����~ 6`'�3�\��^��v�ŇW0��?g�BZ�G��n6�����=���b ��}�p*�p���CJH�W,��7y?<SR�Ǘ��!M�>q��I���2��y�+]����IT1��vM�\>��t <wn(9I�q����I������P�
ܮυ�=I��,W+s,���f��y�h�}ά�5�E���l��%���J�lv-UW�?�����&w��1�+�/!�wC��\��+V��3����B�z�Gd
���q v%��g�b�+�E҇�2<�R��f�d�6ZbE.����Ԍ�2��Ly���m�
�i�{4E�|�j�^�6�y�����P�:�k�㻭�d�!{���t1-�� gw�cxl����%X��{�m�N_��+8Y�v]/߆�s�ߡ[���y$s��
�|e�+�_�(It��^H-:�א��1��s
���c���J��Doh]��3����snTr�;~%p:+�,��Ң����� ���ab*�t��7�\�"�pOJt���UCy�V	
�ѤM���-��?ǟzj���v�^�Zٴ��#/���	���w7�3QS���fhBغ'U۪���ǆ���ܹm��{�7]�5���R�k��%]�p�P������a�5�_b�:��g�_5_xA��C��6�#׫�L�r^�Sm��6dfG�$��$yAz�Ư��T�����;7KҘH�\�n��~-K�8�u��m����&GA�`��
`<lq͕X��
��z�!����b�<t�vF����t���/�ٞP,/�뢷�V�N��>&ު����p�}���#�V�y`Td{��w�!�9��۞"�^�G}�":i��W��|j��B���5�]c��&�&�}��H�X�~�p�������4�95G|g�,�����}�":
I�1����L�G��B瑬g�^}�Yw=R
��[��!��#N���E9.3z7FqC9I�}��?V���v-���p��뷞_�!�|��l\C�S�a��?���B�"CL�/
���э��Z�D�S��kz�'7�b�m��WST`Q��X��|���?tu4���o�(��g��O|BAY��G�J�#l��Q�FV��l��Q'ks��������8t�%���M��'7�-,��
��0sr�"�0d�9��W�ބ�9����J5�e2�������%���2T|�y䤯��o��5�E���;o�	�҃�	�bfO�5𑿪�~.��J�-�]��01�����Y�c���M����hWIm-k�U�����v{O%��h	36���U"�'�}��f��XK���/����ݥE�&�>��p8�M��s��fG��*���`��=,̨�l��N�=(m����+�ǳǁ�"���� r](����F]M'9c�~\C>o��c��<|m��p,4��$-�(�4~|3N�x��/>P�-��Z�X?�i��o[�����?%+d�E�Fߺ��QU�U�O���¹2}F��PN��
�̆�rl߄5㗮A���9=i4�D��5�u?Q�M�q)��8�v"}�Y�Q�,Gg���3 ��&Z����h��j��)��ɱ�6[�&ab�g���qj�0^��w�3��P��];P~ĭx�yh� �Xw�p��s�����'�,!.���Mi�0���a!J�ݨ�{����▇����d�F��Y��b���<Q�n��d��_9�0w�0�0	ge6'�S��?)C<��v�MB�m���U�!o�a�ş�r�����JaZ�<n��W��.��PbS{���}��Lt���f���M����{��x��8w�8
>6��a��������v 06l�s�(���}<�A7���� �!�fm" ��٢|���v(#��S݋g��Ū��P~���g ��jP�My@6�� �������Z����=���������@t���9�ؗ����4����&�j͟�=�ޯ�޺���5l�"�K�����[��G?H��b܆�R7u9��
ml���'c'��yC�_��
���,O��S��M�m��ES7�C�Fe�g	X���aᒠ!ʫ[�w]��cx�pMM��; L��U�n�������-"�V�i�	�����J�1)�k�m��P�k���y-)�<	Q��J��2I�Go�.|�&lL���sd͘.�TQ>�vk��)}_�#���o�F��p�0���z���ioTW�3SL�<�Po�� �O�[��� h�|�,��� ��0�⃒tY�S��V��uEA�|��2nG4���e��&�pXZ��YsE��*�)��ѳ��k1ha%�3�L+I52�c@(a�Uނg���-ȹ�a��t]��\6�(li0I�1Ԓ�̑�f�1����T�75>j�.�]��Hj����=k]j��U�'ѵ���kG�%��������f���ǚڛ{���T�ݰVЌcۮcC��^3��a��e
�]�"	�s4'�� ���}g�!��W��������\�ވ4긶/�=�D���S��n�����W�>�i���_�O��v��G�0�hef<-eP���f��9
��m�ei�3q�����Č��F��Ǎ*j�Fs�"�ʵ�fRRpt���suyhX�b�p��^�C`Ef䢀�O̿�G��P����h���3/��s�pA��c��oFT\Twl��ȍ���n�U�TϢ��X}���~�p�+��Q�n�8z��b�&��>뎵~��5�Qz�ؽi!���������UҶ��őe'`���e�����wAe���4�sU��"��Hu�vV����ineɪcC9oʍ\o��v�8�I;8��y�(|��4\��kHN/�)�S���T�n0B�c:�R�X���.�'o"�]VM.!N
?a�\t��� v��-y�7Y���D����Lg��]�dh�~XQ?��2�������ߓ#�F�T�h����nm�ZwAUr@p�'�����N��q��+�;@��wLcc{��@��W8�/��^Q�����d�z]'\��2���pؒ��W�8.�A��2i9R�d!lW�=o0b����q�SBf���/3N�V%����Q]�Ɗ�t;& ���?������a��e����S�� � ��D`(�l[bWm��~r�E!%-9eh���g!@~lŔjE��j�Y�����Gz����L���d
�bO^�o_�x���Z���}�$�Z���Ъ��ԍ�x���Xv�߿5ڰ�N��bKM��ش��TB����!K�P��`�� �?��\׀��M�n�!c�^�ͳ�ƌ=�9�9S�9a?�[�Q7�6��z�ف��LB���DN�RA=@���\�����(���BS�3��N��<��ǎ������&�y��zY6k�%b���FX($A�%	j��N���s�V��;�f�L@\_.��ަ!>(՞45QJ�rɻ
�s��QD�é��k�P/0Q?�����Gd0���x���)|�]�d��Ǥ�+xp���B╋6rk�c}��I�|��1���QT��,�/�H_R�83�Q�}�J-��bW1�RGen��!�[Cu����H*�&XL}�ե�mqÂ~X�O���jE<�߳t�̛l��������x�u���k.�g�'-�i�hy/���5d8'j4�z���G����t&���Y����ϊs���f۹gҌ��ܡ���(1}<t�$�(�BE������|�b���:��L�
HNO7l* �W?%i�,��H0��w��"]�I��R�[ߍt���,ɵ�����st����_l�M�����Gs�t<}���e�����.4X�p, X��~.��A�Cv��6�E�����OoYX��̨+Ѝ��K���`9�3���8�XސH�?t����r����nnՙ\�N��
�ͩl�H�o3���k	%kJ �dS��q����$�+#��l.��� r�I�4��d�<J�"���Ԑ��kY|[�XB{�FH ؈���Ƚ:�>��_q��YSI�LU�����u�+ʜ�	�{�s�]����d� �S��,�����$���B�u���t��~��5(�Y�OW�ː ��O��֭`�L��~%˻�}��ͱ>E�J��mm���!m�B�� )���X���0~�g�U=�EǞ;m��ܤ���2�?�9�*��=�`o$���\m�=�񇥓���һ����8��hp�/s`D+���rKsi��٨!��Fek�@�Ш͎� Z�
tά��R�XCD�*���Q�\�R�Ć���5�V�|�`.���ݦG�\ ��w�z��q���� g� l�g��M+n($�0(Lذ��F�*rm���T3,!?���F�bx)`�#��#]�>�r��q�k�ُ�Ǘ�SFrA�"��������Nkqa,��9�M�g75���I(��Z����I~�7$��nw�M�ݏ�]�)�������7����Z�yY���ʮD�2�%�ʿ���_�Vb��<��.2����PD�m����f�p?��+��v���;����m[�.K3�ɰZ���n�� ̰:�W���&M�|H��$��Zւ�v(64F�����W��,�g%b�}2 {��������?A��k��Y�M1FD9�`!�u��M��w�^�gHo(ګ�闰�P)~�=�,����6���J���e몠@B��C_���dj9��>'L�J�#f7��rSmy�@��������e�����K��NC#G��w�
��Ü�y
ɫڦ\Pέ8����U�� �l��0��{��Nb�N"̿
7bѻ�!���^����M�R�9bvqM��w���ra��W~��4r�������^2cZ6o1�ж�X�d]~W�:!ga^R�Ɖ&��� �=�i����w���4�B�E�h�=�B|���]���]�f=vᇆg?\��Z��K�M#ML1�?�m���W�59GFӚES�s�C��z�E�@7�P�+;�����}��^�w�-��l?�k]�)u���1/PM6!C�&<�d:gA�!�!����C����͎�;s���͈? ��,1!k��������H���Lb�,���r4(�25/��ʓ;erЧ����5�}�|η;�5�r�[�yN醘���� $@�-д���<[���F�^�qk�t{`_	A��=����;A.��?���7������Q����饪}��~��s9\h\!k5�^��W��Oܪ����	Б��͙��\g>�N���27�yǄ{�\�N�p���?Li��!.�;��B�A�ە�m25�HV����y�T
�X���`�
?|J����់�y�����. �-\�1�y ;ǖ(�P���jWl�홼՜��ǅ�Lґ�%��tu�����d��_&���v��s�|��B!��:*��;��+�c����SvJR�%s�����1�~n�������@�	;i����7:���Ϊ�w�=���Wg Ja#��:�%�<��p�K�<8oO��E�0z�J�.2Y�#OqM�s]�o	?롽qA���j�Kh�hDf:�Ƀ�	��������Ej��z�����u�2�O`<�"�,dS�]F�}֣u��_=_~��&�������z^��k���
ttC���U�r�o�¡�7�y��F���{���!<�w
��I�����p�V�V�|������ӄ��Y7ō+���r�7޳�)�������rr���p[��p� �%k�&,j��fZ��3�@��3A������agOy��_�7�������{%���=v 託��*���V�Al��*B�{eU[��x�i \ߦL�X�]V42T���C;��e:J �F���M5˽7m�B�>����9�_���)v��yH���C�c�gsWb��a��I�a�~JY�k��jh#���k���#��*�d�0���XP�U���zÒ���k�7�w� �m��(�?]�#���z@z�FCW�r:j��)y̨}A���B�m�Y��n�-9]�����՗q0{p�)��5���v3�W�����:T�m.�G��_��^o�'�a>EF?a��J�̩��D=Z�z��y���׼bŰ̷��b(8ݒ~���h}_�iK�֎�9�"F�mi��@?խة������HΩ��� �ä�6�х9v�x�w�G�~�=�#�h�s9PM��r��Ǯ
��⏸���]u77�B��Ǔ�W���c(���4e���Y����Z<�B������ԟ�n��-�d��pU
ǰ�`�=��|/pa�%RB��eu�+�~cS� �l�p�B��Ɖۤ�s��Ԇp�E�xVC���C�j^l�,�;Ǖ��1�	�mm}|��& �d�$�2Qh��EZ�f�y������m�S����,�ɵFz���Mx����D�۫Ւm�n�(������DPj��>��	�ۉJu\��>@�3�S�5w���8�b}w�5�Ձ�
 ���?�`�ɆNg�2��`�z $BP]!�9ԅ���F$O)��V%��y��"�\R��� ��`PŹE���g1�c������3�Nd�̦��3\ߩ���d	��:S�%��ؓ���k������ׯ:�3��>{�7��v�Zo �Q�-��r1�~u�B��g��w�Y�vni���\�P]i��|OFt�]�cȪ`xl�}J�Dr�9�����4��5)u��T�g꧅��m����7���S���f�m�s��B���<j�����xd����d�vN -�/��Z�{6V��#��L��gM�$��_������8��v��T&26qx�����a��q���YG#|�X��Q3.� �9��3��*5�Q��z�#���K�ŘS������(�@�̚�l>�'����,����3�\/��XHj��������0���:���0�+48��K��l/�O	�i�FS�2�C�LG�����OT?��l|̾�����ڏ���K�D����5
���ѡPKI�:��jm䌪���������ӔC{�T>�j�[e3����|�=ڍY��H�.�oH�"�i7y�&pd`R���T��-T-v�yF�9���Ta���v"�'����`�瓴OܔMݳ>p�}�}�Xd���j��h�I���{��d��.��Z��0`w�,�C�2L-��n�"����d*׵i�T�/g�Y�a|{�@�]�^��I��ð����3�X�E����[�C${�}�ق�̓%�[0��Y8^T��jgV�p2�s&58ש�:#9�h���KÐaQ���4�Jh�+���mAV�Q���jZ���<W���>�ӯ�фu���p�tС��<yC��4�T��o-�g�}���	�[�U�KĴ/	G?���������)8��ѓM|�B�wݪ>Yr��K�Q+F��p&�����?!gэ���õֱ��/�ʠ���=�>����#5}! 	@A����N-c��"-�t���Gjݵ�y֧�����1$����n�]lbu�Y�����g!V�'�X�2����-ë�:�����!vE�4$=�3,�'�(W\���|
��^�v E��k2TC��1�S6�.�=�_lc��NS��_���t�m5��T�L,`!�jh�XNk��7��3���n��/&��뷙;F��&�4���r�_� �;��]�ɀu�<|M������"�Nq���v���*e�f&7.�[��}���(~���ǧF�Έ�`�Ox+�����Tm�з#��Jj`�UnC�,�c���}i�F�\��k���$r	,*�:������y��09+��?7�N�1�d+ٹ��i�t��ܘJ@�[O��jUd(�Vn�B8/��)0BW��$ߎ�����%i�p�m9i>ӭ�yc"�n�#Nq�oGP�R}�D&���~��w0�-ЧLI����S�������)͜��9���-Qn	3im[\-N���o2�t�,To�> ��#~18���G�Q���N��Ly�	��9ȷn\=w��VD=[N_*U�*dR��|��q(�h �,�
�ߵ[K<;L��f��-��#)�$��DTF��n-2�7j[%���Hpq��k%��LCL�6z]�]/���R��\e,��h�D�hȜ��w����ͦ���6.���nb�G~��5ɉ��`y:E���R,�+Uc����*ar#����R�p?<�(hjD���T2�����VQ
tB߭��_��M����#�j�j�����4e�K�@�sÀo�"D��'v��=d����y���4���^՗�?�ZF��ۋ6�w��'f��hT���^6/����v�h�ȥQH�Ӏ0����~t׈=.,K*�F(���W#���_������(��beS��l�;�5�=�6�;R�D3�j1�:���_E&�2��s�|ے|G�I�A1~�zZ88kML���7E�ʚ���z��I꿽���T {��N�侩Z���P��3�ݸ�w���q��{]碖Z8�Z\1k��c�ڹ$^���E�����J���Lf9ƞ���Y}An���98 aV��y��a� {d�� )H���,?ڥ+$��#_���JklBq����-"i��
fM�̓)�)Y	���\OJj��NR���)�)��;�P���y]�@�~D�7C�E�V3�eAS�G=���b�L�[n�'��L�K_��*?���$��'��*ʳ_�4zI�՗ۛ�2�~�F�4/YD��U��![��T
l�R1Y�7���M��e��.�{�+�������-��0Y�ڮM�(q��+�9z��LN�X�~
��J�P�];�����..���?�ݰ�ʈ�<�`f��ܬ���`%�9p��z�a�5a0����1x� �&���V�1A�	:�����$L݂ԁ�	���J�n	�80��s��pNK��	��=�Z�`�w9$9,��k�9)��-���u�Y1�|U�7���w����X��6�:5|4���})̕�ԙZ}��N�w/���r��#�Z��Ŝg��*�����Qn�~x���EA�h�[���� 5����n�����0��%:�n�}��7K�_@i��
�j�
�a�����*��/�"�k��ݖ�AC�'��ݒ'��S�&j�)����Y7zi��>�6����G1�#��j{ϵ�b�+���"��窬�jyh�(�y��N�f��h��{���M���h��p�K�\��Ax�ȋV�t�g"��皎E��}�`���d�T��[��L:��A�U����%ⵢ����g�f5�'�G��`�P�ny����x�ivmY�Z�z\#33�F����WVv�h�[��9j�2~uL�4�k���Ph ��jRp���.[O�%����J~�0'˞�:쭢a�����#ާ{Pڐ�W,�|:�cK��0k��������z������X !����}�v�5-p0���U��O�k(&m���Zd<��|�-����� �v����`��E���m/T�fe8�q8P}�Gd���������q�u���B#;ox��l���iםm��@��;i�撩=�	e��Ȱ���+�Z)�ɇ���U�>R��F���pW*m�^�Yb�ة�� 7�D��D�-��}�q�	ux����m
��`#�o��� D��EM$dlN>G��%/���B�˂��o������9��o��:(6���v.H(�K)^�tVd{�Ak��03���nf@u�Y��UI�P��)'!��rrV��6�a�еD��T���K`k�k��ZQ���Ǡ�!�\�l��*�/`���]5���;�*���� �v"g.L��` $�v��'T?�*twss9sW���B�V/f��¨��3u�.�!���r3IO��&��V5�`�<��E�$Ɂ�����{�ҕ�
w���Ti��:2�
�x�"
�k����r�[&g��D���ɹ�rv�^[���o�QB[[��w�
��j)����eх��C��|�����l�����:s�hǵ�RKσ�`����?|��^7��@��ϲV]L�S�A�.,?:�t����fȫ(Wg�D�l��_��h0�e��ߋ���H]���|����Mb��0�R�Z
�<��:(�d�H&�0"M�^�Әē$vcȽw�`h��2B��3���^Y��G�>%C�jnp(d.��Y+<�����5�fG���C�XT��{�Z�q�A��)UA�G�)gE�J:��G\��Gfdl!��)]���0�m�w�ޚ�iFϳ�;f��%��w7o��:�)4a����lB��B���Lbc"�����&kFh08��wvM2��!& G��Acu�v���|A�Z�23Mf�����k��1�H|�ق�~/� ��bQR�k�����2�0��'��ߴ(]�b� �tn�#,E�s�2N����=��"�H�k=@E�c7�ɐ���r��ݛ�Qf�h3�]g��w�S20���Z��2�L��b+e�-��j�Sɛ�oB�僄��&8¥`�,Č�7
N�<no�]Ό:��oͼgr��j�<�}��6���E��3�㷋����ޥ;�hǔ5�r�O&X�m0c�d������\n�DS/�F 8/]��T��;��n]r���=�2hE���Z}�hI�b��Q��_#�[>���c���M��l���:�a�;�9٩�̽q&>����G]�f��1ʯ�@LJ܌�k��
*��� $'�����~VKӒ�s`Lhyt#�1�v�ϜQ�j�?X�����T����割l����E������--Nq��1w�?�������1)�W�4ҹW�ۈ�إ�Օ��CO�|��g�M�$�?0^G4��c!8����4LnM���~�qv��ׇMf(ψ�Ug l���^�C"��a�LE���R����p)���6G?�R{5:p���-�h�n }%<
B��Z�.�8i�O�y��@�2�v�Ȇ����{G.ཧ�U��~�l}A��P�w�p��ֲP�n�s@�5JfٜE�?����W�����3��>��e�_3ڔ�:|Z�[�S�ƻQNh8J	�Ju��S]"ϳ<��D"C(;`��ot};���5�@ϛ4�Y�E����_�4���j?� g�`$/�Ѭ�ia��1����_P�O��$�y�Mq��SR2�z�O� J�5�?z^'w��F
���oنv�����������=�K�s� R{��f��>#k C���5v��1�ي=D�26�\�nx� ]��'�R4 �,[�y����D�}rk۱[`�����k�$�![$�3����-�Exi[��Yv�����p"�R���h$�#\.&�3�? ������3�e���pk����g�n��R���D�����Q�莱���d[��:|���.��g�0)"���&��+�	���3���O�d���f�)��4B���A>�l�qny�oΒJtu 4� ��%�Y&���6��/|��-x;	�y ��
�� �3�'l��c�:�l���t��6Y�,��+��-Jű������K*������D\���]�ҽ�,�غG�.AS��)D�yB1!?Qc4�3�r�[��v�5r��ς�2�Z���$��?ey�'[v��;f0��GD@xY�&��94�c_�⇱�l����e ���#��q	%mihrbMiK���1��rC������YpE�*�Ta]�$�]�;%\��n����4��e=g�mc ��$�_ se)�#ҽ��V�@���J!:�nJ#���ep�NW�Ɇ>-�R���&e���E�X�sH��e�͉�^� س�X�P��S�ֆH������n<)Z��n�A6�r��i�(�:��!�;�699N͊�TLaa�	+���h�j�H/ͺ�?�NA�q1 ����*�d>�El����8H����������S0���m��O3��0xON@8��ah��B�$tvC����e��D�i�#���G�:7>K�����_�͜Q� ��K�v�@p��93�brH	2�9�e�Jl;��d�R�
�;\BB�F|"1D��xk�PS�E}�m0���	~�TO��@ϥƱ��c;���9���3�s�I�t[3D_��Se>*Uom������س��rI
q�Z�}
0�ʣ��"�t]�K1�)"�v�-��;����� ��>�n�D�wm^���(.�j��P�[Ob�8��E�����
�����������\�s��Eٳa�>��C�#�¡�jĿ�����`�"q�ܵ�;>|�,�_T�b��ހ�He\r�ۉ�^�":��(���ð����������¢π��-�GO~f���<�sB��n�@J���J��v߈h��F>L�xM� D�qy����Y������y�8�%~��*Z���1�6BA�o�Z33x�%:vEj����&�R�kP��B>�//� v���S��>��+ה��v�Ig[��q6��rx����y@ҟ���^��3��s_鿐���3�(����^��\	hS���IzYe�(�`�J�f��o�v�Q|�#��|���]&!D���?���޲�-�7�k��Wd�	��9�Yf�y#�q��cB���OX3˛�C��aT:n	��m�$Y�b}����3uf;���!��������i�1݋Gl���l��> X����@��ɻ�A0ʦ�Lx�{��������uu�85�nǐƝ�D��H����kZ� �n�qxi��4�)�5�F6#���h�<~~�H�/��L�H���1��L\��a������K���Q2�0I� � =���TK'lOݭ�.��N�M@��Q7���^���'��흸��W��J������ޒNlhۯI��������	����9#�������� �w��d�dΑI�V�G|��b�Ǔ�~���MW*X�:���$k��P��c�e�4�A�qD��`�X��Vl�<V��c�B��ﲬJ=��w)]��V�&!r�va�-	ͫ��,:&��-o!{�{��	ϐC��X#v���K)@��g����\��+��U�d���ƙ�[�؉�c�I���fX&�+1�%z��\3�uA�����C4������LV@?.]ʢ����`�-l�C����TͲ��8�>������V ��E`[&d� 4���I�3��`2i'��H�!q�^3&�e�r+���
���Q3\�Q@�g�v*��!4~,��۴�r!����0�hI8S��"���L�J=J��<��'��c���8��H%
�ں}��4O��*8ɆFF��5����q|�0�y����>�@U'��|9��"��R-�ܭ����vu�E���$�4}t��<<�F��ҋ����c�GS�`ý�D�&_����6�1�h��E��F��+� �U��£�ϲE�?������*x"|�0����Y��X4��(�k��p�t
����$eioPt���:~��_���I�>�a���j㶱�`��R�3����V�}��B���|������t��p�`����|��<��l(U`L�1�����	'HmK��
\ߒ���^>�4��_<P�ߙ�j�M�=�7�z���稂������T>6����w�U�Sڵ��*�Gz	�a�/)��Ľ�w��V�;��:2����V�%�R�a�������zċ�����64�"ٓ]�X}{�i���Sil'?��Х���h<&���0���/N�a;��Oh_�wB��NN�u;Q.���6�E{�����*q�tW���`��JJ�}�Gh��O����&�tH�YD��@^R�rP�� ��1��o&4SqAfD5Y��=$Ym\s��DX��I A�>n@�<�7���4�Jf'oE��d�)��q�����Գ�T&���ʔ}����߃[�<|yߥ?�k�c�n.�t�c*��ʖ*�4��^�����,��8����gF���U�w�MF������U*�k!��B��=f@>p��8��5�&���*rγ�HǟH���::4�xHȶ4��o� ���5��Nk ��c���@���+�γ����U0�\k�I@x���I5)����7	����Y��4�{E�[��6ӌl͂�D3p�ڸS�Ub�xt�ü@���'�!3�[�^ ݇���ʘɱ�E��9ë�@�Q�3�����4�;�v��p��)d�K~��6�N���$��d�M���{���	d�ːt�DW����dt�p+(}q_��^�ԞgH)���E�pg�o��NT�����Ƿ&�II"X!�t����I��C����@?���B��H�&�&�$ʲݏpE�6P}�Ɨ�6��� � m�ܭ��nMFW��#��o��C�I����o��ʵ5�_�;*&P0k����ZV��ȹy�9v������R;E:��<#��v5�L���)6_In�m������B��(x�ĵX��q��U��JR�L�G�S.J`{�m�-�r��g��HOJ҇U.��u!�E_�Wz(oĽcI{X�u�dw�U`��χժj]�P)��L?v>���؀h�29��q��v�<r��ң'e�y��+NY��VO�]+�����^y���T�Wv1��ek�Tr�UK�I/7D?�����u5�Y�����+N�1�3_|@���7�
�~����v��'ؾυ����w���]wT�ut���P�'5ǈL�V���_:�T�7>�?������<*�ݵnӽ`J��f��-�e�jC$kMvVrO����;�V#���~/�+�ɪS$�Ad�VT��.�����$��G�?�M��m!� �ɠ��v��ҩ_���;�l)Cx4��>�.jH��ː�b������ͤi� � 	b��4��s4���^��審����ؑ������w9Y{�F'̒S�k�O��2����ik����ɸ�����!�z��C��?ߚ�=��a��� Ԟ��臑����Jv����X(E'�B�+v�!��3��k+d=^N�=3��vLXi��9~�
z E�N�ٗEl�ǥc
ip�#�4�}ڰjч���i�A���1
���#9�dt�]
c�CԀy����Gˏ��'�M��"*λ\�*�U&ʈ�KvO�]:I���z�	Ì��%����?Od:�����c*�d�/�
��\2-3�Rb�/�d���M��b��/m���6!��P��,����u-�o4I��|�K�Q�"wB S��ۃ�"=�N��O���q$we�&$p��&K_��+�w
����:�]a����MCQ4��@�8�c�c�f)k�0ٶ�~�� #X��ͦ�3Y�6;>�L��2yu=zZ�8GH����騣��l�3�x�wQ�Wa����L��}$D�#>��*���r�t{��$8|W�Z]a�e!���zt(�q7�@X�G`����]�����A�C��?x%��ْe�h�eL�!��I�eDJ���׽��t�dj+O@b��#_�K���4CuY�m1[���E�k)$��u���}C��v�Z��G��P��MlH_�;�n�%���9��n��7Tn9���s|�0����+V�����}/3��������v*P:ǔ* Z-a������?\�y<��[�=w�'&�O�t����/�"[J����C��1��xj�h����.M�GƜ���$i��@-��	�.ݏ��PBw��mv�V1�t�*�A�Vr��[J��g������� y��:��M�p�w��c%��(�
ާK�z�ߌ�Z�W�����)���%�Ҁ�]IR��s��N'�P�"n���Kj���"�l4`<�2������Z�aW�N�#(���
��!�D�j�������}$�[�[����,X���_����Pp��
k�aeB-A ���C�����0��|�6�I�����N�d��gO�d�_?U���mJ3�y��2�6��+�&�{�~�i��A]�.5�\bЙ}�}T���Z��զ��j��]8	#%�t9ƒ��<�;O3a�'l�߻Nx;���N��,���0���c�HXJvO�<5�)�.�[ص	���dɈ`�ܐ�f�ud���@ ��[��B!��5�gO��bG?<PX#4�ϫy�⼬B���������ލ��G���o%���?5̸���+�0D53Hw��K�E<O��6���9�ˮ�mG?�� .>�-{����?L�T���sS� 7�Ηi��U⍻#fF|�����k�Y�.�.X���<�Q�'y\�Vw�?��Ө	bp�,an�2���6f}Q?n�D����z�Z�^�V�9�9#�҈�j�Ȼ�QG,(Tδ�b�Yqs���Y\����R��0F����
�9�|�7���һ�[ͱ��y'^p�)2e.��Q9��RM�L�t��u�[���b��k�1g����ɬ'	�V6K�"�nܾ�=k��2�'|}�JI��)���X��'j��s7�&�.�|aٜ� �[�}�(�;/f1�#ɧ����a��ُvSȩ�ʙ�{ӭJ��F��/pI��#N��>~]Ý{[�5�^��w0{Jm��i����
��[d?�iZ\e����0�v�l�����f)>O�v�����
�����X�e0|	?Np��� {�*�%
��;�c%0�Yf�&�%�ݞ����5���W����էl�)�4*	\�	�i�^�w]�b1����u
|��!��^��[ݯ���'�Qe�=De��[U�a�&��Y�L�V/���tf��S�����Ⱦoٞ���X�����n�QnhO�nJqs�� �_'��?�T⊴?t�g('�
��2�{��^<��zc♡b�_uI��&�MUSf�����ҍש����qX�y���^{~��$q�6���	5��Ō<..٢k{�d��A0�o5%4ǳ��T�o�wu;�rQ>Z�OaV���X��EHD|�N+�N����)���9�#�9xv�;���**t+C��x����)�Jp��������o�m��v��EVZb嚞V��+ѡ�ݨߚ�bR>��=Q�����ۜ�4��7>#/Y���}�=2]u��朸�:�v�;h2����~bz=	���}���J��.�[S��)�p���v;?��pG���n��Ԗ�%���_H��n����T���~�+�Y+"�F?��rN����]N�_lz�߬	Oo�1's8BS�c��5R��3�Y��N���io����c��A/P'�xHE~4bp�5A(K:���h¸G�L��H����B��Z�7+��?3�^�S���r�:�S_<�_�U4m�n�ɣG�Q�z�����	Yu�h��8�(�J&�<�bi~��8�Ww��p-�z6_��4�~�6��4�(Pw��o喭�
j�Dk��g�Kl�	�or�0r�R@��2�k)[���ճYOՃ[�<\ t�jr8�x~e~j�ʂeYM�����P-mh�YB�D٬HߞlB���T�61��L��ڦ^"��h+C#�ߋY����CC�ڵd%W����J��v1���g�zH�Hl�,�X`q�j6`N��i�SjY�	=H�P?KFf�|���I~_-�L��yza|}�ƍК�]D�.�wu4�\���:���%�K8�D@����N�~��p�WB)�G�	(�[Ee��b�k�7�S9�P��\�+��rd�`Ə�YU��h��Ec�_��ʃ�D�1��ɧ���#�}0YI`�G��kh�>��;��d��P[9��#)B+-wrn�G}�'�nnC{��ǿ�.I��zE��v�/���OkFP�&�j�� ��v��ؘ�����>����.�x��!=���y�L<tp�k|N��^�հ���5z�Bm��*E�����O�d�i��Qᄬ2A�4�p���s��j�ypd7���ͯ �t �ޝ���LP��˥���n���5���#6����+�jn҃dL�8L��ZD�k�^��%{�eh�LQ��'� �.�3m�P֋,��K����8ww#�T��2L�}(:=�q��H�=W�<S`�d?�ËVjk�J�hn�ޫ�1�,jy6�}�r�#;_Ye|�ǧ�
�b,��� G�����al~�zf
&��ki�����(���P���YR�:^	���W����܌�?��=�R����J.R��OT��<�-V]�ֽĜ�I�����e,�^�V�g���A+yP+w�U��ո&����Ǝk,�׫"z��u�0 �+����2�S@��	�ܶ�t�ׂ^�I#�L�h|!��L66�;ھbެ��eOsۃɬ��H��(��%\�kM9r�*�U���	�~��7!�5��"�^_��̍5�t�k&�d�B�������J�vᲓ)=��l�jC��V�H66}�V��d� Q%��=���P�13�s���E�"��Va6G��W�[Q����s�9�Q(n�Z�`0}�Ir�\���p�C����Z$N�� �&/������2BO����q�P߇��a�h�gtM��n�Oa�s<�eX�m_H�����//���j�}��’.9{R%~Vk[��6��$+
�R��\���tC�Ō�.u�����OV[����x·�@N���ʦʰ��(�������e�(*(������ʀ�-����$!~*inl:�F������}���KP�NK?���v��!ٰ�R9Ns�M�^�B²+���K.+���tǐ��H͈Jr�S's�����pg3vP��>�~G?-1wS���N7<����9�kP���c���������;�bww����w�_��WW4v����	O���?���un5S�|2Ů( �ג��$�F��i���"�G�u��`}N��잽x(UH&��߆��|�u�K:ͦΑ�zS��ZbsN�p�f�mR&�T�ʟ��%�a�v���	 ѐUK�+�x%�wJ]A��B��}G���s ��7^�X���s8�_�}�CS���JY��͂F��^�@�
9= ����Z��m�	!�kxo��.�^^��-UoYl�3/K{�~���;��$D�����	 Q^�c�_\�V.�?/�J��d�^jg��bٌK=1��!��ɯ�̴��*$E�(����f�THˢ#�P^�����?.�}������9��6y9~Xd��G[�[8����U��M�ƕ/FӀ5��}��z�K "ҵ���2:n\�Rg��ڂ{�h�z�)��������u��T�Mj��	i) �[�����;O������hSu!�l��͉zv)�����p}���6��z����2�z�����v=)�w�1X��61d��/cC �i#��� ��D����A�n �ď8R;9y����߄�Wh4�R=zܾ���v�-�v���iYw:�m
TF�H
�[�&��Pq����g�x����pө���ڼ<9BP��,yhS���)���3�@���}�}Fvn�x٣���l�lnr͉�xj�w͒�fۊҖhbU��j,a�����1YQ�����tb`?lF���f�ƕQMI�;��?�����R�Z���0�+�0��MH��R�x�Q�p�t��j��3�*wQ�	�C�q!����B>��F���0۫�5*&��*��Yd�;?�-�&�y��f뒜�����A[�+��Hkq��<Ql<7D/%���-u�gB��&^���Ǣ��I�q���=ʽ{��r����Υ�5Y=� 9f��2���hC�^�i[m�ݟa�+8)4y"��k�9u,��Ї���+-;�2��&I�[��2�F�}Bw"f*cYH�R� v�[�m�v�q2Pjˏ�^!�NM5�`מ/�t��#��Q |%LG��媩R@+�d�J�(y���1�R��j��>�Y�M)թ�B`���I�(��&�f���f0$o�
Ȕ�g8Y1�\lnb�z�{aܖ�����>0�2'0��>HK�����R�ߥ0��r��=h_��\8~�g��0*�������UcU˟��eڦ5Hb5�	����>���hᏨ�K��F��#��+����YXZ&�j����ő����x�g]Yܤ,:h�g�I��&�Sﭒ�ܡ$��_�u���| ���T�燒�5��/�1��=S�v�2x���W1��*u{�1�\ƫ�3q����>��8���jg{q��dz�=���^��i}�e$�E;;�y[i����aK� bG|n�7�Ly���	�0=�v.��r�+�9dW���� �N�m�kT�F�P�W�q1:�L��W\piL��\�X����Б��s%w,J��׾C��ҧ�bR�������3pKㅓ�ӱ��H��R ���=񫨔�7N�8�G�y~�d�����?l���Bzi��*l�A�	�b]�NvN7��
���qm�������s2�NH����0�wK{@�Q�� �Iݭ�&�m:<!�����N��a�v�zJ�Q�]W���@�\�C�9�����mxc4�:��g7��m@Cú�C�$+��T#b�Y��ã�O<k���n�h��iai�������k�2'*��I�q���V2_��3T�u��>�d+L�+�C}�^�%�$7��a��"<�h}�D������+�S����3.������p;�1���*�(�T*W��k��@w��v���~�����2�_X�\��W" �M(p��>b|��z�g���8݂���UU!S}x_���}eT��9T�}�/�QJ����/�W=>(����	��@9�L���	*Q�%���bz u=����9�!\~�"Z����W��u�2��ƿ��/#�d�X*�,Kx��r�F�5#ݲu�5(Us,)�T����9h�Pm���5>
��p��"�TE���f�����K�i9�H�o������$b�`��}�F���KC�?�8�b����q��OS��Q5�c�g���3a\�\�P�K6⳷�������U�j?a�����R�W������"�(m��Z�P$�$4fwbQ�?N=b
F�
12N����W�r�>�%�<�vk�6bzJ�2����6�?1�*��{ �j�Dk|Qν�����`-�r~����c�l���ep���(pR�c��9�a��l /��$������8ӡo���Q�`}T=��fA:�
��ÆU���b�#�f/���y.�<{�{�[�;l�vt�]dzD/j�o���@"y@�*;h���SN6э������F�}�ɵ�y���Z�?˝�1�:#{O%��_���k'���t��s]��㥒�o��>�x���]#K�F:T�͔0y��=��|�Ff���+��<bJ
���Q����X	w6 Hbk�YE/��(����;Λœ!�v=����B���
I��?��\>�8��>nK�}�G,���W Q�`��d>6�cf�N	��h������Z93���ٳ�}�s�~}�X�� ��S�����a+ �GV
k|-����`z�@���q���Y�����1�GP 3��u�gǻ?uV� `����Ě�
������腖^M3 ΋�0��c���\
|zj&�/��?_-�N7:V�: �d\���8k䪠|w��\w����+Jf��}�=x@ vhf�9sZ�
�2o��J��:�4y�aH�zMC��i��k�A:����涷�NYH��Λh�	���Bb��+��_p�X
��l�b~ϓ����dh�|�P@�A(�_!赽�!t�w<�1���t�f��M���$��Ӛ�'���)j���Y�7Xg�˄�b�+rw�%�a9�)m^D �aʚ���Juֱ��y?3\q��p|���8q�����*����JV����w�W���$�ad��0? ���o,G%gb��q������(�Q���5��TD�����Gu�TJ���Vlb��� ����9V�Ws�%����AQ�`��=����t�xUϿRsz��PP�j���^�����5_��V��8�
<O�	�"�����0Z��2���� �����s^�y\�x&�_����΢ׂŶ����k{6�њ��x59�g5��X1Jq��NXw�J�z�Va�?o�9dH4u�f��:�"q��!�?��9!������y����Z��pP�PbT��Q��L����I�8���,�a���ǢE�q�l^n0�Ld �w�O���l��3���2:rή9��h�S���t|$�?g�OBa\p'�(�������4*�W0�.��N �csae��R�E����E�LRߛ������p�B��Q�trB;���Ҕ���k�J�ήy;����b7��L˽�1>�^���OqE�T{į�7��KCM�9qȩP��Ο��U�Վ�'��ܾ��nԨ{t�_Ξ7&���
A������T�@x�%
�~A������5ENaIa�� ��_73wcB(@!�fd��D�����E�~˴�ڷP����n�ad���J]�d��r��Uw�l�u�8��C�W*�ѫ�$N��L�U�$�C�@̧x�R��_,���GI�_l�7ee�j��
[(���_���`��D����	u�a��U6�+�&������InvԻFi�ц�-���D��_Db�&&�2��I�~4��@�aW~�m��N�\Y��D�)������4(��5MRe�D�0Ζ��?�t�g���w�z�X�`��Bn�?ʟ��H���ĽŢV���{Fb���G.�iI;�� ��`D&�k�ы����m�f`U�j��ȇMJK;Ŵr��nPRj�yZuq�,���#ܕ]��@B.԰�lQ�-X���;��^٧�,��\"Z�Z�C�i4������>U��d��<ٽ�{�U\���%�����@H�7�@9���޴�ǽ\�7ۈ��f�گ(e:�8&)�%ᄶ��u>1�u&�9\��O�fnБN��NSഔڦ�]v�i�d����O��9��d�xl�WB��/#mmr�g�]��Β���*�mnL(�P[���c��p��'1iP���Nٖ��֊
y�R����H���h9:�ޯ<4[g3�)����}��#�Q��$��C�7�[���P��ul�\���"PL©<!̥�?9g�P�����#��W�P�l�]iZ�f�	 ,��j�)�x�2�i�b��<\ٱLN^�����P�����$����@�\�S�@>�O;+�'�d<f����:���^���O�S��.��� �%𧜶����q;�F��PE�X�٠�����z�)�R�;A����

J+�S �٭�<��Z���B?�	 ?�XPm�$[$��$y�XB0z�z�p�
|���> �p����ko�k��Ҽ������L�����QS�-ɉ���y,�b9i>�1�o�u����^}�N��j�g5ZA�2C�sWs�T?����zN��5�˰��r+�As�O���Y#I��w˷��#8k����Mp��Kğ<�E������[be�Yk��
|Y�D��P%�pt|�LFL�4�q���p0x'�G*�g�c��1��֠N������[9n�'� �݇V"cy"�A5�q����c�����WhX �iÚ�*�0�2�o��D02�`�$+����k����>]�_P��lWn�Yp�I�U|�Lz���Pq%��=�$	���c؍Rrs$t��O�}!i��ؿE_�;� ��ځ�<}j�M����OP�1�T�6�_����WC�,��ݒICp�X�Ku�þ���{�5��r���9)t���i���Q_m*ihmc�^���xi�7���^�↻+��� ����d����X�&vjo��p���F�g��J��:P��?S�<(���j����M��S�TI�bzP^�@���e��zT���`,�ߵ��nw�ܹt���|�� A7�[��ek�&F<�����%�q8��}�����g�܆�:� Ǣ|�g�~"�(S'�"U�]���\�LF�jg��?Uo��פyg;+V#6
ب�&�D8��s8�C#ؾ�
'@O��|F�{��Ö���z��A����9�01?���.u��e��[�njL�ũ2$�*��昖a_��<�1��qA����!N[���c+���V5�~�tT�
)凙+�[;R���������S@��AW
��,�/Q�ζ'��6��g�Dg�J,)����Bʱ!��1���葐d���#�X�W��kȱ6�:�7mJ!�x0"�� @OwiԔU���h�����gf�ɧf�8��ax��(�ʧ��ޏ����x������⮓A�Uija��I��^%�?��I��JÅ�00ɮ�Z�G�;�����ڹ��.�{��n.��	c��s���a9f��:.�zd�4}o�a��NIp,˂z1�z�'����i�!ޮV(�2����[l�l���{��ӧ�s1��SC"������]7TCxi��k�*���R�3H�o��K� �'�^�I�����3R��z�?"����l[4ۿ���/���ݏ�d�/���U���2X�f� C�y��.���=&�n�)\'��w��$���1�|�z��=���gċ�er��"?�,�l�e�=��}#_�W@��MHsGrj��菅%}���i'���d}ԯp�j����{�&!�MD�u)or٨J!��l�:�n�%���0mD��S0tm�����W禼��5���*Md��G�	?JQ2>�-�4\p�H[^
�a��w�l1�{��57wEt����<Ew��t����H������q�0>	Z�\q��2J+�b��Ad�7�Ŝ�+*�_a��ot��A�R�IhR����j	���֋U0����b�v"��9������� �Ɏ���?�"M�q���IJ�x�\�F@n�CqPZџ���#�o�N_�t�.�@h�͞�T�	�Z�w��U���Z��?*�Zzs'�M����n��\
Ϩ-��3@�"���5sv�����F��|w��q��P
6�<�_W�/^حC�Zł�&YG�k���0�4IL#=v�\�x��˂�N&���FI��h�란q�\�D.�%���>O���WF�(�/�ĬQ�IU�$�jxR�{�
��o�P�����q�=��Q�?�����̴����%Y&�kb<)���M�u?A��ޞ�}A�RAx�[�A�$L���aƶ��E��zy���ڨA�	��h��_���0qKKz�>�-<����E�.��t�0ڈxz����`�W��dlO�=%#p��Ց�PzP�z-jz"S�G����mk%��*�4���` �x�<��f��L��i�C�LL���W�E*�n�>o��)��Uoh�Gk~���[�魦6N{�+�T��RPU��.&��+�`	le�XY��͸6���B^��N�s�h`̬~�]�X��|6�K�q�޵�#�%�V��{'��_��w��AN���x���M.���!���W������Z`� -2�%ht�%N�������a�l�4����<��6�>G �	��X2CE�6�97����B0%��(��r�B(�!�e��w�أ^��;�m��es�ң ��ZYh9��bU��f��P��� JM�p��i��a��͊�B$@�k/A���z�?��7:�D�R�?4����@(af�)@�Ny�NL�X �����u rnC����v?T����`��m��8 �E������P�|�|�.��=���
��|���ry�ԑ�~=������Iߵ�TL��vD��+=��1�l�P�{*�o&�R$����8�}�1mVz�|���}�%�V����s�*W7gd(�Uü�X��p����ېl��-��b���Rd����:'�zN�I��O�ZE�o�z�'?��J�\n�v�����V,�s"����	���r-�̮�q�*z�����Pa����kp���Թ$}��/�!��ok ���+a��/&�d��&����k�Z�0�N��^��N�m�Jc�w�Hz�līgȢ_ӭ���v��*c��t~~W2��|(��j�\涆5 ��1�8N��g1�sv��_ �#޷��Uu#��^���jkl�,L��=?J�t�~���$A]V�A�����a�]�]�n��e�@��zĖ��'S�v����9�:�	�٣��k�
��|ue�W���k���_�!�+ތb^�$�8�>��ʝ�I�*x�П��c}�`[�t:�DI��p�P����Md�s@MR�)��m8������M���`��3��l��x��� gR`G}��ֶz$��ץ
��̺�������hp��$(��"w���j��Z�����^�(��<�z63�&�L�+y������6��i��Z��I����tn���􉑷b���;M��1�bFY3� &�c��ʐ�hC��G�&CH7��D��e�b\����|�eoh�FY	�]����+z�|�UB���H���\O�U�
[�Y����Y�����L�B����)U�O�����X��%��A@Y���a	����!мm΅NO�!�U"��s���ҵ�T�?� \.|E��/�=�OC?q"��ɀ���ǽ�k�Dv�>�N��]a\U��Y��WQU����kD����y:	W�"���4_	���-�Ѓ8��&ZfmB𴷜��������
���c��;Ֆ�T�Y���z�yBz�u��"Z���=JI>V3�!�[t�0�Ra��'�����{�B���q�ٸ�q�6zܡ�;��Mڗ5�)z�{t���|� E���>�A��+��t_X�����V��A�v�s:�y	J�&9��{�B���m�5�
�j�=��4�Z���p�G�]��1�}M�8�����?LdO��.U�&~���%��^GFd���lg�?�"k��[VV��K�~��QUK2���b=�C¡C��x4CTy0$�87�R'Z����3�P�T��^�Y�����L���s���T����ÇE(S�}Hn�|�@�Pc
�њN�˨���rcQ/����?!��ԡ%e��C�=6�g)0p7��O8�b7�2�EB2��I�.+2����]�U/YQrGc�;R��$� �*tg���d	*�F��<1[;y��P�.8aـSC��[[�l�E���7t>�.���-C����9蒒��R�O�6I��Ȍ�"�!~�N	7jCo�Ь��
��)�#��p�~N�Im�W�����	)��>-s�1݉�.w�쌵���9��@A�^m���t��ia�C!h��%��0� ��.��y��Sh�����c>���:Ŭ%��:)K}{�-lPF�$�6�5��  7�л�����W���%���u^B��HqBu�^[�=d��({�*Y�On�<x��W�g���z�:81f�g�����_�����xZ�{��=�0��E"����S��-� �kQ��ńs��e���N���}i�b.\�L�9�D���M<��^�i˯�wyF�+��C���9�1�b���S�5�>�1��`��1�r�I�������.��dld�
}/?B��a뷣�!��JtqwF�uC,`?�HC�E�}*�Z(�bq��j{��<q�.���p^����MVa`�!���~��~��<�+�a��\�~�%�tJ�}7��+_
��۫�oƛ	{NR:B��o�q4���U���B�>z�҂y<�7�
�'X�~�c�֥��Ӵ���tk�D}͘�r������U��&�\�c�5�3ǹN���Ǣ@�B��0���h
w� P�^�f b���"��ĭ��9�������x	:V
�aa�����"_��}��C��Ճ^����a���t��4%�_����BL5� )���<���BFc~yX���}-��=�o`��c���۸2jk�c���rY�)��G�w"�V�3�2�g���~�=yK��4��Ip��O�y&���@8�r�B�>��y�x[*����-��0y��#]<���	�TD��zf��Q�9�Óe@V,L��R+�@z\��^����5v�aN�~\��>��a���2����p�^��t���D�0�X��ٲ�_�҈p;��\ԃv@��:sƞ^1��O�C���d}u��d���y�T�#n"�#w�|���7�6|b�$���:�;[
�sc���M�T��jw�l��y�2p�K���5F\���lp�!���%_�Q��G���b�y�{�,q,H��Hi�bc[�s�{�|�e��G���>E��(5���E�T�J��\��L��4�+.m�Y2ḵߖv7�xO={r�%�Bù� ����;�HU�]�뺎CC*�ޡ��WAR���Q}�n��'�K�qf�mmP ��5L�وB���&�πI(7������K�ׄ��Ȕ���I�v~B�W��M�c�z]���Яm�}�X�����$�N~�۴�K�.Cl�PK�"{���.xxC9& V~F�$�ZehZ��7x�� ��P�[ˁaE����������5��� ����YWf6I��`,�we��x���@vE����	:�4��c�S��#�����-�u@�Z0���deI�8� �m�>���Lzz�%G�v@��I���`5�[b��3*@g�����	Bscc�А��{x�� ;�����O��.����V3"�l�*���y�򁹑gSor�|�Q���Sf�t�ҴE��\&���߳/��a】��N�Ϗ?��<N������G�.�S��0DZ-P��lcw���WV�9��0��8�?�p�̃;��`"�_i�}��KSl���駗m��[Y�XDa��Hܟ4�@^z��!g ��Bي�^0�D�A6�M; @:��,���Q�8�=�(\��-��Ǜ�C�3kyim� :˳��5 �X!`�2�з�Tn�Wf�JhQ�pw�4{li+����<C�G�y�=_���'e��fCЋ��hմD��eZBѱh?����(�R��y�-�wq�%=�()�2K�#7z���(���e�1�Pn��=���j9��0����ji��ʅ�b���=��'ƪ�P��ᕟ�MDj�x%�G����!_$u�T)LS�$�R�0�T�(�჉����{���D��oش8�,ʷa���qW�ɬ<p@.Q�/��J}�@�m�y���M���콭~�2f�4�"�_�J������Vsz�q�;��^�>�(R���o���¼Ü������TE�����բ�v�u&$*���e�%��R�!+4Uϵsq�4��щ�&����Z,�އP^��^���pegKgu�ټ%��{�E�v�w�^*U���l�BF�[L�n%��v�0���'��ٸ�������|Ǫ��ܑB͜�W��S�m���&n��`�Sb�C6�:��{������&���b,.la�e8�4 B�W�8�:�xl��.�>�Ji��U;����.���Qy��AY�_��O�6��j4�f����X�Ǿ=_�&�����@lYT.6<k�Vz7�I����?�;��/�2b\{��e"Z��m���0Т���mc�ē���-Xlk�Ǿv_��!Z���"k�X-������9�N�!�/�ѽ}�O���ZvNw�+ۧ������ݶ%=��h��c�Gy(����<&)5��D	�p�њ�'��L�!�i��Z��SiG�9�s#ɵ����0�]<YTi�r�5�J���W�C(�hG27:F�'y��5r���*^�ׄ/Ӵ�c�~&�S�!(��x��t��𵯿d�~�(4ݳ��$����}�������K)�V�ۻg�/h+���'�ӈ�.v�ы��g͔����J�۟ì��Q�G�c^5�aN��&�p��v��Q���-E=^�ڝ�4M;��u�y<�`8x=zmޤ�`(uiP�szmH�K�N��U�����_K2��_�9�� 춞���$��>���#x�4�f�'�gع�S
�wUe�ҭ�I�o�3hx!,*�`x�nb��3�����vפ��<���(�X��#
�7�K�c�-Dg$A�dd�����Է[��C�<�D�S���S��^p��j٢.�u�x��ַ�C�~y6J�^�2�ֺ'�r'4�pF��qk�\�bШ��� ��Q8�"e7��l_"��dz���"�K��79�VKĻe+Dn-&[|�"܎�����/rme�s�
Xh��8�*}">Rd�޵*�W����T?7��'�u�N�  g�����<�j���,m�ք�)E���ip��D��r��T���%M���_QXl�z�Mҭ��*��e� ����W� Q�����|~�I40�]����I��h������ճ��<cFQw�
f;�А��L�e[��OՍ�h��loh$����
�q�N5��ѿc;2 ����|-�G���W� H���%�u~E� ��T�h���%E��x#���֫��m���ڭ�Fio����h�@���K���?�ܻ|�S��B������RL�_3ڴ�w�7ɞ���?�WI���������@H���M��<��p1��{�&L��k6����'���|&7�?Y5W�<�1��A`���ȳ�H�<�\�%ԯ :����$�p��onb�n7�hQ�=s= a��`.$���Y�b�5��э�z� ��K�|�Y9V���Ϯ�����0:Fhn��&M���b�r�������FKCd, ���=@���5s9�;�["W;UX�~j��/�A}�n:�h;!�oL�ֳ�A��%��dh
��,�7�R
��l�Y/5�EU	���O��P僫	7t�+3/m�NK���T0Gr�O�Xi-Dzݯ�x��.���4m��
�g�E���9�ȉ6$0��1�5�;�R�r��߰��p��LgTj���\�X�gH�ga��F �����$������F���{�}'$�#�{�D���-
lKQ���;�Í���T �Yg��ώ��3sIs�U���蓱Ϛ�9��9EvE(�ek�T"�@����H	o��IK',-� 3����W��멕iJ�&/7��pS��-�	��5(\�`���آ�$C�ě��c�wv�@8oBل,�"s������T�����]���n��r�׶�gt���ņ�Y/��
Z��h�6?�\0�6?���wDb���`�'.Q
�O����a$98�¢9b��`�h�̦y������@���Rl�����/4�������u��q�`9����-5H�����i��H1��~��i#��P�	�n%F�څ3�]B]�~�>	h�!8"6R �ҟ�]]�h�`�)���[}Q�/���ӵ&kZ Z��k^�Ж)��\!��Ob�~��}�Kh�xS�N'ԑD n�E�I�G">�Ui�`±��GL���bP�vf���}���3`f�{�壪jzb���2P�A��ң+� ���Ys>�_:�T؟*����!���Ӈ;��P���k�v�(/X�&���Q�ڭ)���jv�q�6��Z���=�I�����1�@�lv"��Z�`\����1���V֫vp��3�O�sC��Wʃ��E��Ӻ�Ԑ�L3l.��=/���������ф� �eq� 4�~��?n?V2.�(
'=�N�H���_�����s~�le�^�AQ{��tu�*8@/��'�'o=}�ǋ_��F����\��	�.et�"N�;��w����Cb�[��/�� .�錛_��Rl1�Led��gU�?`X�r��)&�!\(�H5�B�R�����ԍ���s���Lg�w�ꊠo��џ�s���u#�{;�C��X�md��k��(����taΊ�\�|��ǋs<�� �����-�fS'�2�h��0��aA�t�Pf'
�!+飑���N��Bn	���!k���_�"�Ξ<��!�YzV��4q��)�m���7��g��T94��sK�`1:�������W��nl�Wz�uBB�����p����v�;,ZG��1�O8�Ң�k�0�w lP	����0���O?�|�5��@���S�D�ʟ{��_���9��'h���so���Gy�Ç�!�]����H��]��x%!������9�e<�B|�n�{�Iz��
�Xu7g�;H D?���^��]�>L7����ulăn�r)�c�qȷ�p����r�k�h~�`�۫�z�o�NQu�x5�f�I��//H�Vd�T���_�٩�qM��B�va�Q��SlT�0�*��w	f|)���<���v�c q!r����8���֤��{�B�m>g�>��R���� }
���o���ջk>��x�gi{9|�Ә��v2'����Y��]�KL�/O�f4�lv���)��BB�@ ���Cy@;�:�}Q�tM���w�f���`�K?�+PZ���.������?aC��Ǎ��Fup��T4�;���R����ۘa��"��x'����\bUw��h�KT��SX�6:��]�o�G���L�8�L�>���q����j��աMq���2�1֋����&Nb=`E�����0#Ucޖ����(7$m��w�OIT0�q����6�~iN �+�l?����h#O��a�M+Gݻ�g�D��~�D��d����ȓX���
xh'q���P����JyB�ȧ@��X�2�7��aF�@�����1�Q�.O_��VK��Q�l�˪\���c��M�������JRh�V�д����nt�`6�����#[ˆ$;�.u�ƺ�}R"4ވ�~�F�[�=-[�@x�2�
V�ALA"lC�[���V��s�}���%{�D��U�Fv��3H�g|�l#7�l�b��[v�� �`:�p)E�%׎V,�wr���£��˱v������}Y���T�;U��Lc�"��wz�Iޠঁ����)�_��H�M�䦰��
��?�.�u�c����`�gI~���/(�#�rj��0jM��-h�+B!��~�Gt/i�;����т�6�U�>zU�v,d~�%R.�WO\J�9�V�.'Oc6X�ʦ��CMi�.����+:�3�ݕ-�g	'H_0�AÓ�sD_��9q���#K<*�1�Bˮ�Rx�>f��k0�'�YP鸡N7��Zʉ�}?��9�>ߛ8}�����`�H���V_Ima�&?z�B����'y�d˚V�쫠z�_���/5�BwZ���$��=.�	s��<�/��Łx��aw�l"v��[ �/����$U�.��W�f5BU�����UP֝�6�x�z�o);*S7�0")E,�N}ĸuvR�Ι&؋gO�6�����9#���?4Wά��W���i�� (���
B�����R.>�o�����^�G�i"�� ۞B��}q�M4|4�R��?���q
1�\�����02���ՉY�K{���f������Lʶ^
�'�a͚ݝ�U���>1{O��L��L��d\C͂+M}�k���H1����7�Y�a�6֟~��wxﰲQ\}��Y�c�����"�,�r?����;(cu�O�'��sR�rUL�z�ݐ�I����9��/v9���D�D��쏾�r��']�����#�Q�.W��;�U���Ý�"��}�V��E*kSlE�����DG@�r�6�T��I��"c(\0�2��6"S��x���7��=�ԑ!/�	��R0�3����گ0�3D���{��f�lX�z�|�����|�ףv60� �B���df�aa��A�i�B���lq�r�N�^+��� r�Fx<�k�6���W����ئL`�`���*{F��Μ�)6D�nI:�|���gf���vƻ,	����l����ݧ����n %4�ɋF$
���Y	
 �C���8a��c�T�9���+}��q�W�漐� ��1[�O��|���!�$�P^��ou�#�!��ԧ
Lp���2k@o�vjt,AKi�{0ϥ��p����S���T�/��b
O��l������U��o*[�l�������n��E��ݨ�s*l*��������Z��폻,K�&�-�<�#�G��'�L�s�i��6���o��5��i�G�7hmF@I^�C�f3jJ0=�P�|t'�;���'���=C�ն��r
��0WK�8^����	�	�{`��u+M&@tHm!��ޛ'��ѫňL$mc�T�Mʫ�����Q)���࿟��.�P��X�,~�C�OG2�����RcF79�/]���_G$��\�e6��!�'\�_7�WA|Rzx2�RP\��r|C�>����N/F�l��I�H_�O���V�s"���o�|�*�y��9Tc:wM�2F6���<��.����x?�:�8�(:�o8���Վ��8�-#'�$��h�����j"~��X=l�����������g�.01���d8K�`j��Gj�:���l��i�US�`�'�M�)L��<B_Uz��5�.wH��g��>@�pRs۶��_�6+�'�K�`K'ۉE��g��՝�bb0�@�5�"�P�f��gމL��� }����X�x�'h�!:��gϲxa�H���n0�p�bD덚U����*)y�^T�4�r����t�c�cq��V�����L�ӕw�A�k�ӴЀM!w��Vp��Tu&"x��3�?1�wY��	�P���R��y���Y$�{�T�c��,�+�_�z��0�QC�ʀi�r��[#�k�܅�8�Gʓ��8�z5 ,v�� KCN�f�2t�Ԅ� gس�j!_���o���&����o�c��K�-�8�@)�"��9�� �~�b�lyv��܃�9�ay;Jf��bF��a2�7��ix؃ܼ-x�ZԜ �m�������fv,��J���й�T��8��.mQ�ݻ� ~��#�#��Iㅮ�����	��*�^=z2)_$��S�TF�`�� ]��88�>��֘�����s7� q�c'[dc�D|׃dWj�w����n
UO�ǻH&!���wM?[�r� ��Qk��n� ��!򡃋�Yz@�!Wb�!�Oq�9c��Hi�{�ٟC�FNۿ���@%�K�6 �0-��mX�ͣ�#��y�0B�1ΕL5�ο��4�aT�}��~fp,D�@���#T+~g"�AY����R����ؓZ����L۴��N�L���3m��"�Mb�ʩ��V�S#	�����D"��1B��|sf�����XV���k{ݴ���d\�����Vvům4�>���+���q���7�"ZĘa�P4U�9r��uт���}��{W�4�y��t���fή���x�n�F5���r�]�p׆CD���)��[JEW�Q`�[l��H��z����՝�Yޓ=.~W�ٺ_RJ�F:�+$�:{��3hU%0�{�x�#	��a&q�?vY0w?`��a@U.���$��^�&���i���Q� w�yF�)e5A�<������ڄ���;o�_Qw��'�ލH�]�� �2�Pq�˥O?�3�2�荕$l�F��������U�p'$J�>"�R��e�KB����㯯��&�Y*z�J�
/�6�����5&4��-4�\
~���;�.�J��:<�#���>]���b��Y/Ϛ�$�clv��WP�C�Թ$L�+ˌ�8V�;}�z?��{#���C�Ɠ�+��o�ɚ�~@4y*��W��J� �x��t�<T�.|�cTf�;�m�,�U�����[3;x�0u��"܎x�Ԅ�����)��N���b"�c֤�!Y�-c�TЇ��|G�~o�������g\��^� /I��wOxV�=�Vl��i
xBWT$T}'��y�a�g��f;ӏ3e�5����0�{��ܹ�]�}��.���b[�������/��%�k>c~G�bI �;+���묾��~���w����00o�� ��^�q��
 �xf�./�32'*�n��T����]0Sf�/��<M $z�<�>�;��q>&j}��� 4p-n?�J�w-p�{8�Wv�����k�q��[&}����sgͷ���*���fR,��K�*3�w�.aD�6v*b�JC��A"<��m����%�ة�Ҙ�̥Y�n+��C3�)�>��'��:�\�x& �����|w��^	2Z����"�+��q�:"+����\���|R��9��,G�^�}����Mk�Mx��X&:1p"��I�E�c����R%_J֤.��x���ǵ��'f`O\��J�,�Vz9[g����  AQLg3��_@m�Ȫ)}���
t0�6���¥��t�t��_��e���w���~��U���X��Z� E�B��^��3��*	Ŗ�w��M�C�J��]�r?UFP�GC�x4�H���� B�q�:K���O;U�My���L%p���� n�ιq\S�GL��r�y���_ˀg�ema��,��fq����Ԛo��^�Q���<u1H3~x�KX}�e�dg���+Ė�_ܙ�]��Kg�vmZɮ�Hu�K@6XV��S i�5E;8%�s���fI���u�N���ՌY�'|��:�	u3����l�wX�� �*��@���jnRDQ?#!Y��b51?���e��#V��%2֜'ل��ͳ^���9p*(��ь���l��[���]�aUlDЅ~�ZO�I�TE���`;gW�ߣG��\-?��S7ꎚĲ�>�:�}�ǜ22<����g���p�p<�mU���9D��S��.ł�哭�x]�ƀ4��%��u\�,B�j���;<�0M/��h۲�\>D؛U8Rޑ�DQ&��\q"��FO�8�z�[�-��|3^M��`���{w�5ݶ�"h����2	��T�����m����	&�C��#�Vz�*���X�K盓�q����4��x��`}Z)"���vG�� H)Y[�F�x#Y��,B�t�e���2e|I7�$�R�\��Ж��\�dw�+��bN�
�wk�,�O��p��&e'Imẗd�1J��i����.�EF������XkZ��V�[/zJ01�\˻,ZW���nמ$��32��Ҝ?�~`G�0LRo��˷?��`?�=L�w�d ��NL�(����Ŝ��߾{��JԺ��Czh�\ xm�E��i���M��ʉ�c����|.���w�}@�����]מ���,�k��S[05Y�N�#�&K����oe�����I�b�{ͅr�`K_d7ߊEO�8�a�7��e�O�l�h��C������=��LcJ;�c�.$���Y��00��ӄt�[��jK��f��^oLT͐���s�B�����vS���2N������PҬO�@��>��^�J���vic1�?�♘�$�������pEaֈ�7SQ������"C4C/��o�6�T�1n�n�-?���{n�\ar_�;�<H�b)@\jD�,T���C�όfd�郯�{��[oʑ��R z� r��S�}�oq4ߋ7e����\�C���b>����!��'vv�s�%�ay����O����/�%�����;����u:���'�la���@���dlrժ�������	^s�i[��!
�Y�j��PjЛ�{ImDcm�ھ�4>&� i�A��b�28�����,���"x�
�J���4/�L�5�jtI	�]��w��e�J���sw$�L^�~J<�8��3Cj]C]�-�m�ŅN�J'��8]��1������P�;�e�Sm���p������?˹��!X�� ��J��)D��^~<����Y��5���0jNH�e�h�Ȇ�_ִk���|��/�xl��A�霕��Y������aPPu+�b����8�׶��-�z&�P��}SF���E�8uIrnwi��GA0�D�Q���mbWg�u�LR3�j���euJ��D�D&�������������Ka:[�$NmѺnwq��g�B^㵢'��ǪcXG��Uj% l ,����K��r��"G�*��D�I��G(��D��.�J"�jj��J�D�4����D���U�)��/��W,3��xd@%�Гƕ��Q֘��^V6�:�:�0Lq1^�"��{"�E4�/���X�w�7��A���]�Da�?�-W�t��o������LII;�}�Fs(v^*v��n����U��{�x�/��|�籶�� >F��~P���❽`�^?��J3G���`��9�4���.0�O��jh"�HzI}E��l�jr�c �ԯ�'�MA�e��4�m���\䩧����<�×[rۉc�4*J��I��
fɓ�������z���h�C�w;���~R�j��Q�E��#ٽ,�YS,�I�~P3f�= �Jjﱞ�@�V�02�k$�47�>�D��Q4�x]��{���D���*��git�g	�[Ӥ��������%׿�k'��(}��5 ��'��,�h}\����,�D�4����M�	�`aØ4��W%�v�� IQ��m!����)���E�����N�j��E�Õ=�M��:�{��]vd=�W�[Ւ�
�k�®a����e�ژ����v�������s��P�D�5�h�٦�iZ�6����;)|q�3�=f��-���o�O�_C��9rK[ivy�{N�;��Pro��p+�vR늞D
F��x�mv�bׯ���7��&���(�dϫ� �7EQ�MF:��M�j�!4ӕ)��.�y1$��!w1����m����������2���1ʋ�NU��z�[a����3��z9�l!9��^)�X7�D���A�5�~���K8\!e�2��D��Q�j[���M��J�mN�R��^}^6 7*/�y� ǏFm�1�tZpV��"����V���r؄�; p��;���M�`�����4_��1i"�ښ�4i���{��
������a_���	�:c��c�-Q3��!Q���NG��EO��~��6�05c�W	F�c�}S��A��H8f s%�aXJ�	T�k����8�׿�������[�ik/~*(D%�id�G@�^�¹ƅ�e��T𬽔�۠��r��ǐP��F6
g����՞�4ҹN�$��j�#�����O9��>�H<s��p�v����Sd $T:���D�:�$ث:���dTi��p$N\Q�U�ho�S�t�-�} �.��NM�{�.��(��M*gnUTH�z\�L�z<q6��<� �S����+*;���*}R�cq@m��F���7B�$��l0�Y_L@{��y�|?yd^;��Et��H!�+Ϟ}��o�$�G�H��fK���a��@�v֡c/_���"o�L��1�ע<]��w7�놦p���a��0~!�WL ��z݈A���J�T?���ac�3���J�ZRuy�>]p ��_����4���jI�GzH��)�=M�ݡ�O�K�=�P2��U
�,�/I�Q�fevfk�~�ZQ�Wy�����Z�Y|�P�ZViM�/�t�k����rJ�V(	;�L�E=�ۊ�vZKC��.�?�X��Fjz�Ps�a����rV�D�M5�2gh���$|�O!f���予_۠�A��2͈�Hw���7�%׷�<�'�ӱ{t2=��w���L�qj>z<�ñ
�"�)�o7��φ�9��Â����ߟ�7Oj�i�2��NR��|�S�����.O%��X;�\�/�`�(��DI����R��o1����<��[y�hr)e��=��Ac��k��|�!B�(�̸��A6�l�i�zb]"԰3�vALO�DB���n�i��|WV<�a�;�o�pEY�V'R��j��:� ��6������y�+}�}�g3E!��{�@�����.�����b�Oo_λ�R�O$��O�hy`�k��T�nE�|	ǆv�xi���=��S#��i���أ@�d�=�T��kvgѠB�:���xO����w��)���>fev=Nfp�x�>8Q<��UNtq��T�����i�q��=E�o�d?R�g:m"Q��6�1c8�<�ʮlRO��Z�~�M��8�j�P��]7Q�pG�+�rF�t�e��9$�My�lL�)��FS�WA��<J�[�x
q���'��xQ��Z��6�N��z~��n���b	j[\���i�k�a^Ɓ�{��"&��*̊���vV��~+������N�V����5�0��0�&�R(
&�l#���_S7-C���b�B��ݫ��S���uk����O��ix��ơ8��BM��L�x�e����/�]Y��^VSc�m����lxEҁ���rNDñ�v�i$�)���tM�*����3� w�,�W֌����da�$�z��Db缾�pHK�����kuxzc�W�[�@C��"���:m���{8� �S�署�P��[��0��:�.�����=�:@];�rZ�	������E�߽��T=N@:#Z�4� �w�����B	���6���4����F�H�����!u�|lԸ&�b���!m�K'�����9��ǐ*'�A��7�~ޮG=���.ӹ�ܵ��V?�5�Qg�D>�7Lp�Y��[C���ػh��r	f�Y$�H��'��&K驅��G�F� �V�y\�A)G��Y�"���f�q��(�F��5G�?ۋ�~�l+[��8�D�GH�)�
��L��P����kY���
��xPi�I��Ď�A`��t�&ϸm�/SJҴ�b���r���y�C��6B�l�{t=���"x�o�Z̊E��by\D,U{�-ϔ���hV�|��B%����D-�?�5'ƷHhj��.��kc��8�A���n|�izޅ��'����20���j͝� �e!���2��0�^dۀƇW�>�_R��Jj�HY�̱>.%Rk����ǽ���\�*����ҥ +��|�;����˹3%��r�Xf������������<�2�n�kq�$��F��&��8�ѓTO^��������xVY%��a�?��A#A����|���L�rA(g�`�{ܵ���C�u�Ͷ��KЬ-Z:x��#Ul��+>ۑ�2��M΢�(w�r�*��ӻ�UP����W������:+,W�I��%���c\Y�}(g4��Um\�ߧ���:��zS�56:�t�+Bl�8N�S$=��x�?�+�)���Ѭ����1�vO��D�ir`�gD��6�cYmU�����E��n��q�y��"�� �N�]�Sl�ņ�&�h�1_eW�8�����
�����pyt��)������Շ3{�/)�����?�+����"���3�n|�G�`H=~��G�jA3SA�6�_,�p�^5��2ٲ�"^o��!�^z;+��j[��b�F5��:�!���6��z�GV����K2�
����s#��l��(�ڠ]+j�ե��0RD����:�Fiu�='��ޫJ�ƻ�ȗ���GN�r�"IJ	.1Ȑ��|��}eM�Ksn�ჲ�u@�{���Ϫ�ނQ�+��{ƿK���)Kh�
O�*��z��Vll;�>��q��)V�_�sg�ua#�^e�F,�QGp��a����,D�x�i���0��`]���[�$.*�V���\ϪOw�,j�f4_K�1���̒�߿���㈪"h ���j[�[��w�s������P"�e`j!8�N0k3����kh�M�\�Y�(���S��P̙�U:��h$����tBgE,cۇ4�@x�R�����J�1=aFE��ii��Ѿo�>硓��l�mO�%cI�O{7g��G��_�<�J}$j8��']����Rʳ�X�&@V��k�$�S����	1��V�`z�)�ܷ���7�Ʊ�����H�+�l�r�ᐑ���]֋�4�|<I���'�5�Ҷn6#��q��Ӛ�Q6Fq&��ƹ*U�c'O�e�>j�4O3��٦X((����'w��G�3;�]4>:C�ҫ#���tƁ���R�=2O�^5K�$���{p��d�[~�~<�`x��@�>���/t$I��)��u�zy#}��i����:�,h���4K��Q�'���ڣ��y:�^e_�pQ���{Ԣ�T7�Ľ�'n�O��5�:�8ӏJbv߈���F���tT�MU����� ^��Y�����>����A���A�~Q����s�����V��;Q�;#����^�p��� �[�xx�&�^�l�BCn�
��
*�B�@�^k�J�O�21�N#�����b?���D鑉�""�?-��Է��^�A8�wk����T�֜�/΄ˁ��yAG��y\YlUD�;��nx-c�2'��$��,p��t��Z{V	�E��&\jGd�T�7E��c��|2[cG�����(���'��%����=#Q�>��L�܏(D�+�Li�B;M�4v�P}�~��h[�`|�yD���ۉ�>���O�"@纸7���Ma�EO�V��CJ&�+�R郇��<�"8�����K���I�0�D��$�wH�[����0qj92��(-��&'x��j��.яC�6p�h���L�kBX�{����r�]1�Z�h��̛��]� ���6�w�k�2�����
s����0U�bVB��z S��6#n�Ⱦs�yBMiԪ:�z%W��%,�o��N6�DDo�>�s�4��q�Y�	�eb�l�_q����m���J�2�Ik��!:×��PL���������>�_A�!����C*�-�6i�_�����ȴm5���w��5g\c���StB�̃	���7�OIt���	:jL�3��?)T4qb�(�SΖS32���D��?� ����lZ�hX҉��Ӯ�A��ݖs}��DO�_�ձ4\�1�!|�ݜA/��b���:˰w��Fbŋ@�x4tY�'i�bsEZ�6⣁����*�l ,t����UY���-)��PQ\�����29��Wf�����B�xi����2�O�!FZ#0����I��m�������/[Q2��7!IfM�e�	�LT8�����q�J�`@M�jZ����y��a*f�b�3&ɚ�8|p��4�n���m���AaE{4x`�xψ�zXB��0���i����V�Q�`�8ΐ�QRfИQq���ۤ�:�~ n)������q���������w9�i�"߼��
�~
�,N��S��ۀ��w<�^��S����~:�K y���G�ݰ�G�?䇤�z'�j���>t�I���$�$�����x.^&Y0���<>4�C:>�Y{�wۑ?m#fע�Ya�\_J&)��)�+����^���+�i� H��v����܁,����A�4�A��/�6�����V���o;�Y�g�T��m7�U!ł���t�?_��ƂxX)u�F 0�_C����4�h@�W�����3'9)�W���u@���w`�����id3n�)������}I{�Cݞ}`g#���;'B?�)�+2G� Y�~�5��܊���G>��R����
�ݱ~'OA��j��=>O���\𨟁���p���;�6���=gG���Bxΰ�N<6�ǻX�.m)QJ��A���{�Nv�U��)UR�~���%�ommæ�u����D����uj��i
�۟s��]g��8El.#��w'����VƠUf��X���x��̸b%؇�YM�h�^Z�AK`��L�����>�?ٙe�*,��@�d�٤���D�cRMl{�d�=����$��w�)�>.�؍.�M��%�R;�qR(��v�(X���;�/ΑPjy&��^���O�����a��A
��I�%n&��,���U, 6�_t��˂���*��3"SOe�����%��L/8�py��Q��Kg<{����[ p-�Ƀe*� @p��� �B���@ؒ ��;O�D�V�#P����ԥk�G!cR̀n�-�ݐmR�#4����r�?8e w�(vV�j�\�+ua��/���=R������-�F��v9Df��?�I�j�8�:7�����+={w$^�:�SV���U����N��Ұ����"闖5��u���~tH��q�e[F�Gp��?���П�*DQ�Z��w�JE��"̳����)��a�V��Y*ǫ���c�I
�L���L>��2.��[�i7�K�-�X�]9�­=OoK�0l��n���[^�*B9r�Ls\!�7�^7���Tk 1kE���ە	E"�n�*����DCA$Z�����U�->�uMш�&U�ᰘi%/1� D`��Gp&T�y�Xë}��̨�wx��6�q�-��r"��pa!���K���������X�*������Ci'"5�046:��)Ut�;���|Z=��s�}mn�U��j���䔁�S�01�Qr�E���P}�cu5�����T�5d��L:6'��&��M�x�i��1aWm�۵Zub��8���	�,4J��z&�a}�n
�x�����M�Q�u\EgB*ٳ>g���r�C��e#���q<�J��
>x�0S�m�-�o���'*Q�&\L���	�$����!z�(��c�f�?�ڞ�5�����+�|�8ڹW!�F�����4��\�ٖ�/�E'UMvc�o=�ۤ�&��p�:-v(��T����+U�>H������ʅK��]yT�6QqN��c����� ��M�1���n�hˉ<��2�lx�ِB��u/�pe��iܡ�g�k��%�n�����``<e&��ĺ`w��4��%�EG[o�Ȳ�9]v��|ֻR�US [m5�h�s���]���LEd1��^o�ùO��c2Xp0ל��r7�t�Cy3C����b$Q��������Ặ�np��Z�\GNa��5���u��Jv�����*J"��������^#~�=?oTQ���=����(H~��pஹ5ܷ�g{��P��r�z��ˊL�^e��}}6ڲ���m�]�]$	E�M����侟�&6���CT-#=��,�{�炞���C�NJ5d"�<n&I;("k�j4QC䳿�E��KR�Γ��rw�2Xp�� ��B�%�7�n�0�����,/�r�.�I��ԯF˰��[�k�.O`b0%�o�;��)Ga.W�ўE���M�2����XC`_�L���m w|��1�&���16���S�	fB�܈�D�a3����S��*~<�.�߼z�
i�����DK��|�H�6r����?�]	�<���2x�|�i0��-1T�j�#����U�OﾜM�w�&>6�Y���AΤ��lQ�jn���~Bix]�0LI^�R4�MӠc�E���q�!�g���K`�B0��X� �h&�SU_�^���B�}�SI�{���v��`ר"E�sX�P�3���2�!�4�J�%k�Gל�ܸqDS���֓����-�B���YA�[I�;���&��޳9�+�5�f�.�V<����i��Ȃ������:^=��Y"���N�>���s9�P��[s�	�i3� ^�j�z���Eo%윘�)�V�[M�Bas���.�XmN_�4�W_��IJ'�zU �~j���)��d�,��þ��3���1�P/�tq�f�92J��7�?�����I�3�#%��6��Hb7���ż�0&P�"�?PX��9���K�c�4C�Ο��gԯ�4N>��Q�r���E;q��t����~l�O*G��@��$�����M��;�K�J"bN���.�Sa�,�-�1��4�=V$&v�!�-�$i3ȏ��4[�,� Y�^��BnHF��@�t���׌���Ёg�=�Y�3[꜏�|\���w�%j�>h"��i����`��#��K�i`{�K1��H]<nq�ȠҖ �@Ҭ���5���m���
�#ؔ��e�]�Q@�Z(姆��:C�e��G3��S(�ev�y����ܾb)����z�����g�RZK���ēz��D��4Dbc�4C�9it-/gZ�b�K��E4޺�]�����h�� ��h3_��
c޿��=6V��q
E�b�j��M3��ESX�y��q;�	�ʓ��q�q�s̷ii%u"�(xі��3�-
.��_�K���W���b��(��
���`�A}���n0���?�v�q��#��O��a �K�J�ph�)�r�cO�� u��S�������k#�I-�Q�h#��ܖX�ῳ��{3��_I��5�41�?1�xO��F�`�^d*�T�)�3����X6�0�IF�8�=���:��a�EX�)�Cg�Ā���)��a���!�L}xE�o]F�� �mE���Yp������Cw�8��6�p�}Nҷ�0hs�m�kp�w��ȪJ��# �Q����]�1���L^/����C!�r����s-HeP��Sy_�X�1Q%�h���U�j��$�j۷��(A��H�-��u/�w6���?�<��J����ʹ�^n7n�F�Ξ�_OCj�a��L�.���׬���k���+��m������޻+��{��;���eƩ���h�$"!]T��Vt�ۿֵ��'N��Ю�)�8�"j�?ȬV4�2|��/�<���]�LJ"Q%�V��C�~���FN�J�~�\�pƌ;,Ļo�ׇKh���-&��LG�Hc@G ��ۭ>��IlLy+��|g.�I�ƴ��+��/o�6�D�t��s�{���#
v��pQ(w�i	��u-�%�0����GZ�:�	ec5��������c������TbW�V~�� 	�j�O���A:yv����Ƞް���{��s�򕕊��	�ϖa�Eif֤�);��xƚ0Ӣ��ZW�u�iv��Ι�gu���iL%�zE%��>;�Ci��s��Љ�P����%���~y��>����3n��u�=#"�:�=xM{JGZ:Y<�y�
��WvT0�D:��Z֚���{��$�~7k�n	��n�8!в�،眙:#�<��'��)Rk�^���(���-� @�2����u׭�*Y�Ձ�k���Ӌ��EC�,n!�����:�����0�y�fh틟Ol�$�
���R�bפ� ��C�O���_îU��. a�Kgw�_M��\`�6K8��8�s�`�N���Ylu��sm����Z���>����1�F����Vn]������>�l�}nK����Li�R��ӷ�Ő8|�K�"F޽Ԅ�G���OV�6WO<;:�����*���}��M{s�&��ѾZ�(�N]t5�� ����Y�K�����\YPɬ�3�(b��2�Vut'�v
�%���,9�U�
);sL�"�����_9)�~�oXE�k���5�VG��)�"^0�/R��vfė�.Z��j5�VրV�� #�~�k0٣�����E���;W��`m_�O�3�,�uߎj�f8�q�Bd�8�/8JGnF�+*�g/�xB��F��T-�������M��D���/��a�;m˒1E;a���U�+��!n���Y�劃��#�h�݌rHJ����G����5�Yw����G�@�d�8j��p���C��T�Q��t�M�7q�,��F���O������unr��Mc�b!5�gE݂�\w��;�}D=�:��A�u�>N[��h$��*D�M��L�Uv\a��Ы'Y���U�q�#T��Z.�
���e/��7�v�ץ��I�h&8o]�(g4�Kγ�f�Y_`�q.i� ��4��=ֺ�yuE����ej4�X���l�̤��ԫkOWO���3p�y�u�����ǘ�
)�>��ݎN�P/�̚b�Aڄ�ޤi	7��W��Ͱ	t�9����_Vb�%��4�i-��w�O\!OeJ�l=lĞ�Xy��b��mJE(���s{T�ĥW*�{�%#mUc)`�GD���A��β����^@Bk_���MaYu�T��������"��`c�$&��Z��e�2�
s��ݷ��]��<��NH��Wi�u��w��*����s#|� �Õ�#'ez��z���c1�q��X���S�+��2m�	ϯT��3$�T
��V��
�8�]������;��Kڍ>�1P8�}��-v�K� �6��L�|WH��\�����������ܖ(T����]�
�&$���@�Z�=ΰ�n�Y�Z�#��/ǉ-ԍ��\B��gDS�6�	�H� �	��}f� 1}�E	�ɞ[)�)���YL�6c�I��;���0�ܿ >Ⱥ��i�}xW^E��5��Qs�iA:���:IW!����tC�S�b\db�F����.�m�@����1�^�	&��a���|�����S��S0EV�˦�:�.����¬�겘AI��Rfx�Mb�`낾8����t6�=�"apZ��:���&4h%��W��b���"?��� CWL�t2P���oA�}G������z�����{qW'�!���������/��?�������%T9�ⶀ-�G%b�;�J������-c'ɿQ���FJE|���	��+Fa9��˧�V�ȴ��xuZyL�2sx�L�o��G����|{3&�6�s���Qn�����(坜WH~�eP�-��#;R�s����-g��pa��jT]v��~�ԍZ~58�'M��p~+O�]������R��d�R���ˣ-�,�n�]"�֝`sj�0�7��Q�E�F���7���lƮY�������m��m���!�ŗͯEib�Yn�3��e���Q�z;&g��p禙'o,&����J���q*��X���
�e��v�M�� Ǽ5\��yN�tBd�$~�����}�H��H�B,0��O���z�T8�(�l;hfNc��v��wp`��X��hEcn��pd�y���ϳh{u{�"��*��GQcY��-M2�$��'�Q�P���픉u�$�࣏��I���f�o�Fw�m�|�숋�R�E�^�iA��R�?��J,��@���l��s��o8��N�W�ڿ�g� �@^����#2g�Y%X�v��'E���o�������,m�C1�y�7�L�=t���$B��Ѥ��(�"aa�JuZT�b�?вL��1U7��`�UgN�$�Tߝ
���0H�Х�Ɩ�v�c�8!E���q�8���B�jO/�7p쫏�X���d��]/a�_�Ckfm;
 WPZK��G�e�C];�������12�G1T~Nr�c l��S��bB�d$.u�b��-�*����}Ou�?
ky�46�� �[m�g�����<��z\�Đ}7߯"�B�2��;�i��q&��o���+SWp4J�H����/��t�H�ښ�L�2N���Z���l��)ccE}K�DQ��ؖL�1��Ch`��(IF��׋߯�[�\<�Q[.�Ṉ��q����U�-�hR$�'�����pmY�tg^x�p��[G�qS���P>3�[�S�Oǯ�V�D!^M������f��b��{mLy���l��^��M�����hMD�H�nrP{��ߥªߎEe�V�@��d�A��ʭ��W�I,L�`���|�g���el{E"�Q�}fs���U��'�UA�,���e@����Dyo���bW�Rk��7�"~"h9z˳�j�X\�[��7�3�=g������Rf��.t�|��S�(n��V�	"��Dy9-�E�!�xZ"���b�{�W��{�KA�+�3z��U�s���
�{�1	W4����GL��f�\O�
@d�mr�xlt�įc�!��L���Wg�rIdʀnߩ���.�rtg�@�Ѱ��rf�1�F�ۆ����oK$�ݢR5g��LA��v�@ ��kc�hf��� ��(MB#f<�k���x��ԡ��,���`?��X���Ԇ"�M�<��(4�ʳb6�d磀�q���w�R3��'g
�K Ac����;����qbB�=��f��_����Y\�$��[�0�~��!���p�k�h]�-}zg�Av4�(8\TR�S#+N��\�bo%����b�w?f��Sd�)rQ����/�8Q�&(��_'�k��t�r?Q49+����k���<�d���mse��0��w�1��n�}V�����O)ͳS��|E����R�]��r��S�n:��E�P��'g�_�;�4��wW�uQ��L���a>!'el�(v�A�j���_0������Z�K����7t�;2HKde+�!>�$�bм?�2�"*c�y�,�/�mԮuF�v
�Ӗ��ȏ=k�|�u��l$^�>���� �����H'3d��Ω1����w�焨�æ�5s��GU��W��� �Å�7�r�������Z�)�I��	�j�u�^DG�5MX�z�Gȭ�uK�@�~L)w��#�P�؀�IzDe�y.���';"''���ȉJNa��D�����-�W�nZ:~a���f���&��ˏߣ���i��bU1�km,�h��8L"�"�<�{x>��ٽ����9��)A)�i߈}h4���r0��fVHz߳��L��Q���\p�K���YL	~���o�����;6,C��k
��;6� ��$��À�a$tA�P�����gR!�j�7��~h_N�.��OsMS4�'8iq�g0���������@��]j�Zj�����u]� ����� �ܿ@F����(�Q���=��~UD��P���X[�����>�e�>͇V6�*��c��F�~�Ǝ�1��g�
���*���S�2��ո�����E��s�t ����k��i�o��aFO*|��x�0s�`�",�u;��|̏��`9�Xݩ�8����0��ɩX�T�k�g���5����ɦi�כ��G�v��)C��"�}���s�If�lx���$����?O����,�p�-�H�͟�5��yP�K��s��ER�B��I���n�mb�{�îq_�#��ǳlC[vI�Ru(��1c���Z{�����ev��*Y��tq���`�$�������H�� ���|�t;{#��Iv�.��H�/����ҭ2� Ǆ�Q5N+�¢ک�a[bȮ}�7��
t@��Q��ڝ��$vp�j������$�f\���,BxE��2�JBm����_�|:K�ۿ��kI�Ci���;�фe��bH��r>L�S���U7��!=�|�d�|�!Ŗ/�0-��Ȓ��H{�n-���G���U�)�X��ɺM"��)�
���W��	ym �(�E.���Y�|=�C�����Ŕ��[wLn����s�F,��*���F4��C���U>Ԁ^�i�f����d��,���t�YT6SO(H/��>�t&������4ݱ����"��B�"b's��������.x�ז��E� [���l��t+�86���n��+Ft��7�E�+56(� |`���m�*�;��3C�����c��*;d�s隄f�谁%t���E�Aeӑ��	$�/c��S:�;��z`����y�����-?����zXr��%�I��e��se=�#�vq�6�D�c���v+�72r�T���k,^J/��� ��Xxݤ�8G!,Û$[� T�h��3���w��"�E�}�8஬t�Y��	eT�]�?,��-`X��FB���VB}��X����؉g����{ԧw�P�[��D�ɷ��Y|���||�Ù�ѯɹ�h��"�iZ���Ɨ1 "�ENbl�t8X�Er`G�Mz(��c��(N{���2�����8m��
Oà���{���ŷ��v�E��D4�ܔ�$Y^!�u���g�2X*��d��$���(f&�Ж��d
(`}��UK��l�����A�Ԛ���У J���~�Îl��R��ނ�����P+HC��eC�]N���);�����J�̠pjT��T�̡��Җ������`T�-`*8�ɜ�
B	K�7�_9
�Œn��}����
�K?LsN
F��
<�<p�X4�3r�����D^}@��o��_Fh&B�^qK���$ET
��%��#0;�ts�5��$��I��9������H�-�~���|���M��0�ל�׋�^wd�UyZ�ï���M�]�X�����za3=�@X�N��<�Ҳ�7����o��P���i�,����F� &��Nu�d����$�*
���Ɵ���>���(��|���TPW������gfU�r���F��J,�d!��ؙ�B���&?�S���M�X��w����u�uI�/���[� mi�t�����$�:BrT,��m���`�R��M+���M��Ι��d�n�'*�>vӸ>M�P{<I��@���5�kK{9;�:��?x�
�Ry�d�e�R �g�P�H�R�������NH��@�P^;��u
��O`���]�a��������ӣ ��M�*Hp��˅�,�i��{���Q�d-�N��}����M����q#S��)��mvC�i=��?�W�)zrJ@B<A��S�����[�`9������wN�w�7�/?�E�����5Ɨ69�*�ҨuG�WoC�]T�|>%�Yl8=D�<�&]]����8.��gU%���V 0��A�>���I G ug�o|:��#�&�J&5�a�nQВ-������L�;�nw�E���AKe���������95�6,�>���쳧6���sq�a�{7�^��6k��u�����*��$��$�I �CB�N*$?��<d�Prb�<��K�b�L����c�NHZ�+o�%r#���}{y�>U$-���V��a�lա����`��D@����N>��<I��3�	1�\k����g�� ;yfmf�)|E��\��EJs2ث���_%�qx+G��Od�(l�F���=9�WCDz{W��e����!9p*ی�Q ��c+�z�	�;���"��(��dH�
��8���L���t�n��^
�2�V����y���!���nǦ�&N��.����2#��eّ�sPT�ZSv�1랶��z~��F�}܈z�}2��F�j!�?�y=�Ώai�������ð	φ�}�Z{�����-�����Nj�FjQ�ݯ�$m^5�@L��u�q'թ�&�%D���qة1�PM��"Ċ�ۺH��7!_�6��`8�\�S�c��p��ͳ�ꬅ�8�M����,x�G%�j%�G�y�9F�k��-I�q�`=�a`;㩝/D���+���_bX%!��Q�򽂪�iX�#I��;��\�K�6�!lg���S{a���⦨x:������F�-�X��z��rK�Z�<�g�~Cj���Г����WD��`�-��4�`ipe4lunE3�_�u�0]���5�בB5�0K�#���τ�i\�fڣT�Bŕ�1u:��Fq������d!���&j�bt�&:�
�8�/Kw�p��YK$`!#�qi.�3l�ם:¥ڴ����[q������iF�_��ɭ>X#��Wv1�mfWČ�&�p�Qr.��pq��vA�sX���"Z����4��s��9�p=
��B!5�H�Z@��q�Fg��Ɉ��ÿ�dXp���X%�%K��_yY�~R{��kh�c�{B>���4�1P���2 ����NCy����K��.�P%G6X��Ͷ P��l�f�ը������b�rm^g��\�\_0���;�J�����3wh@���f�ZLXT+#�`ȧ�a ��3�(�<Ũo�|�-����\�*�,�	���0S2�|lJr���ڱ���Ѳ���"�mC�)m� ��a�(��/��aӓ�-.��:��-|�|V"��Ц��r 1���Ԥ�e,A�+��ˢFF�|���E̿?�%/�Z�\1�5OK5��aN�pI药:�T��Nc��'�Ts]]S$���Fs�Cs>��v�0�R%��[��c.V�Y�z�����h����o�C}����&F�^ʒ���o�t��C7��o�E� H����!؊@ڸ�cV43�|��0���1��y��]h,`!�,�0m�P=HZ���pw� �*��k��%K�������#�����ѲGI� �eR�[² �B�_��� -�H���� zhe����g��x��I�3��g�{)�����ojg�rr0F�;���b�o���A�Ef�Y��|f�������0J$�Ƭ��J�7V�>��� o��G������p�n,}mS������5�DQR� z�_Z�3��	��$�A[���ǁϭho��=wʎ�ۜ���n���*Z�V<n=ppP�*�䇉�YVp�O�����Q�A�$����g��$����2��剢�A���k�|����W3�p�NDB��������%��F{I��d�O8Ƶ����ݰ�ж�����GY���[�u�C��*����da�����(��ʛ{�k�-68]Ws	���ojFcA� ���+�$C3�L}���@��j;�����J޾��@y��*E>��&o�,�����x*���E!pc�IKŴ����}�ݩK(^>6�X4%��8v���A6��/E�ܘ�6\ O:M���	�;��Ժ$�r�z�	�Vp��h	��`�
��)��1?�M{h�C怠�hG�`��-֘9���T�7�-#��	���\�{e�+��5¨�Ȧ�+Tϫ�-��5�l���y��]Ԗ�7ϧ�dBd�];ju��P�D�����d��}�*_����{g�����R-�@tې�����>Љ���|f`���r��|�����	Y|��ǟ�?'�d�I Ĕ�fXP�U��PyO�N>��0@誌yY�n\��j.���8���u���ȥ`���/�T٧��L#�JG��A�s{�~�^̻N������}��lf4-�z\�:=G���v60�p�S��I�����X���9��H =�2�����LD@:�rY��!�Ք)8���d�#TRpC�cqٿ�@4�Y�#`�
����Ok�]�(�lgNy�F��4��~��8ӧCAu�c���v�+]C`��x
�`��)5�]��n��h�d8�KHSG�Rb����~��h��J��>;�!F�N%�I��� �)Z��r�k�6}�3����q��q�xu�1����i���Tw��Wl<���%�&�h;+�<�[��d��؃�oC��`��znP�0H.S�� �����e K�y�p��[-�A��E5���p�R
G��q�{����jzg�!Oj�/I�H�cu�Ԃ�x`(����/�
փ)�a��u�#SF �#�k������&$�vM������Exo�����frS�?F�c�wsq�ۣB�ü*�liju���Օ=n8�߆�nT����"u�
-(�@�d�Z��;7�<e38p
���H��]|��ՙ�	�a�? ���or����<U�z,SR�m�K���,[#���N����؇�?2�&�Ng�j�h]�7g�6a��a,X��}��MX7Q��VI������q/��v����z�p��5b�ᤶ�$T�M���1 S���NS/�g�4�m�<�!��g��.i=0�%}ô�A0ۭ�с�߫!�4y&��z��'�ԑ�C���yos�=ߗ��˂��fܞE�Z1S�L`�����|u���� �U�N�x1�/�k���׍Ld�����s����Tŝ��a&��>�^���)�w`�$a
�6~Eiئ֤LP��g���ǅ,I���>L��#�6>m�ʹ�Twm*@����R����Q���T�.�"$Ǽ��Qx��8���{��4���G��q��z�3/���w6��om����M%��W�t��O��Ҁ�y;F
2)��S��`��oUI�K���V���7���������G^r@9s���B�F�hI�)>��3UT�7�-��:�^p�,��@}Ǔ0���bPg��Wy��Ɇ��-��U�k���զN~B�9��<U�F0't�[�T`�1J_��fU	;9�Ǯmb�������J�=��f@#Vv�46-���("ŽZ��3��7���1W�p���^ �:�D!^%��9���k���+�����.f���5Јwcg.;����Ï�.���]5g���1�-�����YpGX(]�.����K��%��Hq�.��\�.���_�F����a-��K�+��������ZΜ���`����Ԅ���5��x�2�����_$��Kܽмf��d̿?q.+��l��������u0ODVz��Xw�wTT�� :��.Cu���Z^��`�����)e)/����������=F�Y�+Հ��@�4K*�3H:�r�4m���&��dܭ��9�4dϐ���ɄP�^q�E����]M3��~/U�۶g
Q����鞁�2(�o���i�1۳����{l_�w��� 9	H44�����Lʰ�+g��I���;h�M�Q[�v�\!}΃x8�2GD������F�f_��`�`���6+��x�o}L�m�oۨ�h`T�pj��ay�9/۰��Ơ��T"�)�?�����teTC���U����p7�:	W��H,Ԉ8���7��-����xt)���"#ZYF��35l5��Ց�\���"�`�Tm�W ���tAwk��~�ȉ��OY$(=ͥM��O4�5[S�G��Z�B���˭�=<�0�"��OI�;;A�`�~QIO<�W5lj�
�+�-2X�^���Ӟ�H���#_��z&m�!�V�3�+\~{����d�fpBs���s�ܝK��|T�+�6=g�d|mՔ�x �8`d7��pǛ�������W�H犱nu�,�hW��+&�8�@���:ʜ�r���1(�C�����1�V�W��&���ɒ!ҽY�;ޞa�4��e|9���v����v0P�KR��T6���ު�{��|jX9���EO�=-��Bf v�E>��CZ�/!����4���� m��=���[�ף�E���O���j�ˑ�e�8\ՠ>ExV����IU[i�5��J$��lݾ�[wp�ǁ?d�h��Mm���Z�]SjK�6&#�˻��}�DUV��z��޺�Kq�S\����K#ADDuU�H7�Ԩ��#)�~�����,��+am]ħ�9z�|�5y�>ˊ^7â�oKo\�IG�$��^��p�G�/��p��1k�H���U���"md��"�$�"/�Z5/�ߤ�z\wۂ�l����K�q���l�/��
X�	A���}�q�#��ְ6Ec�y樇��ډ�{N�#��~��*���cWK����t}	zj%�Zk�Asߴ[�T���0���T2�͆���ٱ��`L}xC3ե,�P�������N�ҟ��C�#0�#_���tU4�4�
����gl��|�:���qJ@Ɏ�'�I=�t`@$йb2���9�/�%X������y�%9MY�U�p������q�!��UO��ac��v"jj�N���ߥaK�F��O־����q�5~;P!�jg�Qnb;~J4��d%�
�u+��g�v���Y�[!撾�r�n����03�{w�M�瓛��;	�,q́�m_���#8��9ߢ�6���K�L�7l�h��c�X5�����O�-�'z�4��C���H�ϱ�+�A��B?F�t�K�����5?bZ����_/E��{|�!��9�pι�t�	����i��*�X�.�3���;��C_�MSK>�;���7�[�U,�s0�OŰm�2���:Tf]�V$��DZ͌[�.+�+'%Z�I���q���b�3�+��[Cw������]|�/g+J����=��ab\
He�B=����EgT��E�ͤ�h4�FY�}LuKd�O�fi�rk�MW�ML��g4h�H1CV�M�����clƛ�uƞ�K~zQ�%LF�1�=�b�k>vl�K5�E5j-�ᘄ/ g7Đ��6��H

���?;)a�u,�} `u��	h��:��UJ�z�
?��ɤa�*{D���/<�=,���S�Ƒ��I����&�5c@*��"��>˨����<[A������Я����󯪐�C�i~�j�x<�̷����1�'�Qr��Dn8��B�~�j��J�l��� 8�`m�Zv8��������'��X�W�L6)
d�-/cJz��&�<�_��5�8M�Q�o�3� ]���	Y�c�&�}�8�I��y�_�L3�e�0���8��6E�9i����n��k;��j��N?�X2+�J>0�9��N��2��drzK�I�,�R)��<��{��o����.>�玙��V�7�9ȴ_|�%7C�/
ͽ�r��%�$�v7oU����YRW #dm�l��P�{>+�A�����KK�	�xd�C4`)¯���p�1~�p��E�n�)��S����韛��j=�i��eb�<H�wO	c�d����H�����n?����^A,2��>��r*�}Ҭ�6RJ<� i����msU��2���<I�>9x4����������ڧݴ:F#2{�Pgq/����c���PN�~Am�qm�����a�����u�_�xDc�c'3ks;?1,��P-odQA�e��*n��3�x����`�&��Eԁ����P�)�|�<�J6��|���4E9�ώ~[Ⳉ��� /w��WL�b3�#o��4�j0�e�g
_ :�}���-O�cP>�Ճ?����ˢ�c4�S~݁����5��ܣ�y.���w&�O�n1���֗��Ĺ���aE@��|�;ް2d?�)fӔK.V�Ř/X���s/M���H���<R;I�'���&6HUy��/�?f�~ /)�پt� �����5W����+��ޭP���IA���k���?�u�;�SM#n��^H-l��c��ǅ:�̢}-k�*�%��Pq�8g��[O#"�%��w�k�#b'ۺB�ժ�ճ�`��l�X|q�~/���p����7��QPl]C8TD�H�������.@0<d|T��a��&���mD�}���b���{6��Y"���,����Ke
MEl�_�Iê��Պ"ڶ���p�q"�b��ߠ\"���6d�4rz`�����g:�������K�12X[��PL�؜��n���TRM�\���$�� 
c�h��m��	���6�W��ⳬ����Ņ�O&���m�JlZXjG����_kʨ�K�������A\�(����j��TI�ꣻ�R���0�~���{g6�i��Ԟ�����ߨ}-Ƕ�v?g�a�P���Y��̢]B�%]�>���--&p�R!P�&���뒣`󻋰�aC%�O6#B��Zg�>{�=E,��H_���tGǪ���w�%���iv��@�8�&|����;MϺ�|7��:�P�Q2#����Dm����-��BÓ�u�07%g	pR-?�
��f([T*�6�>;dɖ��(@r�qjYzK�����{so/o���<C�/�%--�T�D����cHY�c�P���&vRF�,nS*@�wV
�q�䚮>6C��n����<�Z�z-��QΙ(S�pn�e����ޗ�qؿ�-@��DZj�v�܄/\�2�ɒnk����=�ɮ���bCFz���ό��3�W���	�x�d@I&W����w^������M4u�)��d�����=�X�c�\�=
0����v�aKכƅX��Lj��<P\s&j�n�B\w0�O��q�4_4ڒ�х���ț����ACV��0މ�,��#W�s<sEG�ִg��v�o�Y�5I�E7����Zo���_�`�#=4�KU��:��rX�q�f���V��ۇϐDj�<e�ە��3&����o��aS�EI�Ԭ��h���d�;@3�aA�KLw�Л�J�,V@�Q���xB̿��yo9Ϫ��2F�i�Y��̹$���H<��e�j�"ٖ?I�i+͆��NТ���ga��N��Ҵ��6��c(�����V�4J�����д/Dw�w5�3>����GU�R�إ��=�j��6a��L:��Q���Rr�ʘ1�,�d�6��,���}ҿ��@N*�֭m���l���D�ݻY�Ml�f#� r�DqT�����R�\��u
�j#�n��<����4
۹"�B���(���a%������^�:P8S�AߚU�-P�H��ڀ�7�e�� �ژp�iN����\�#��J�*�%��*Vm ��#�����7Р&�<���C����f� S6��&i=|���o�{i��M�9 ���>�!K�A>>��mP�,�F���?��VW�����M��ǈ0?�W�W2-�fū;��+�A�g���B^��!;�c�,{f��r�wW�8=$�zx�ƞ����T8�ۣ�5�Aer8������F��X�����dk�?|g�˄a�!J��ĩ�#��-��D9MF�Z�<�����ő�~N���e��l�W�LL��W�%��P���q{�⏼���H���9C�WC��uѓ)z6�%E%��״���F>�$�`>���������qmz�S�LY�9 �K���j�g:���j:}�u���+�J�����Q��,}l���/蚛����G=��#�����v��'�9����u}��HM����+V�&�z�g��^W��O�*f�	�\eHt^gڨ�� }`.C!�k N�\蝢r�������so�������~yZ���USW�H�va �w��Q��/t�x��ަL�m�hQ���ů���n
��.rY(�P[(�=c�{m����@���b�-�;B_�:h����u9�*HH'N��3����kR�ym(� �J�K��������鴬��:�������u�D�VOI����6�dً͐KT�og��T^г��{�;��x����Q�����C5�X(��]�g?���U㡵��`J<�7sr�7�m)1'L�k7��̼�|���LaYSq	�D�6�)t��P����a$j�������ґ���w�c�B8T�Q�W����Hx_�$u���tE�Z����\�uM�N9#�������{̄�a�5S�P�D����4�ڣ�2��o��ͪ���S}l[
	��+���#��ip6��3Rs^�׺�?�i.���O�**&.~�nw��Y�ME��	C-�\��Zv.�m/*1} �E;�Z�"��/��?�i�N�(������pԉ9�ٹ�E�6�*9��8gy�+�e삁�*��}�#���\j�����#v�*��Λ�r2�y�i��Cf;ѴA2Jt��]z�.���P�Qk1�]� 9�Lu�W|4�����g@��e�X��;���������X��Ȝ�iхS�)�eD��-�y2B}�[yg�{ж�u��k!/��cف����H�Щ��xq�}�"[�qF޸����E���a��3#���[��`�jA�;̤J0)��_<G�ЛL=g�u.��Q�^���"���9e�d{`uc.��Mx�,i'��_7�8�	�(zׄ�����oH���m��j�Z���6����+y�@`𾭻T�p#����9!����y?a����ۍ��,M��V7	{oS��_�aB@:pf��R,I�W`2aBG`M�Z������,�)���(5���e�W��G�vq�	���^z� Ά����SW�n&G��� �w�(� �����P���+��H�*�l�ʩTef7OC�2#_\����6�M��B��o�R;]b��/@dz5˖d���R܁���6����b(����^�3��W�����H�p6���O��B�owY�3gq��}N�>���[ �|v��:��mP�1Gđg�:f�>��,=K�Z��b��p��a_aT:'�E��[��4��GaX������k5��=|[���U�g���H]x�~�SAQ��&G/ad��n�i�e>�O�g�eU�G�r.cf(<��m�ѳ����N{%�W�L$*`qȹ��WG[Z��%�hť�Mm<�lz\흗E{�`u��/�1�]��S�F|�b6{ORV�(��#�%#p�(j�W!,��]2r��4���MO�<}Xit���X�w�^��������3`5O��޴�H�gg��>�� y�x�PXsa��8�]s�!B��L(���T�ߴ�6�}i�}�-ϳ��?�'qU��:�?5�.z��	�ug���^����V�s ��VoB\T � �$IcHŶ��=T��-��q�Z�P�94�~��{eab��2󓔺�E#�$�����GV��c��zzG��n�&�GS��:\s~�I6���3S/3|92����|�*҆�g~��-�g$7�(�,�eE�@r���ANt��%��La���>� ���ä�/�ݯ�ڣ�7
*6��sw�Z��j4/h�����>��M�N+�B!3�Ng����v�۬�V������<��A}��|@!�q�w�ׁx@�m��Ν:����o�τ��?��t?kK2�<!��B.���?�X� ��1�9{��Y-�ф!��D��쒷+�;J�#y3��@|�G������3�	��F#w"P\�7��[8@�,}��G�4�������!������aݝSv Gj���PO-�\#�W��S
T����m�˙��q@��
����*�t�|^!>�a��ܟ��!���U���G3(�z��֝(Tz5���i��>K�*�S�1�c�ƃڵQ�x�s��ޝ���bJ��q��`�Ǧ��*��uҜi}��{��`�"Q���ڒQ��(sܶ]��C�Wru;f���>�E��`�ٔ �
�ة�S��B�F�c���x�o��;I�w5Y��{u�>�+N`�|Vi�o���Gf��b) ��AsѕX�Yj`�4"|�N�5B0�a!F�<+T!�TW2E�=�58ҩ�Ϗ++�]b�kP��O�qev��)V�H�ob1��\�^�D�)R<籚}g
�Fd���A��K� ��;���R���cč�咧����~%>��=\q�ioM*Pf�f�Ч_׬�hd��I	�_�t���m#��.�.	�NM>|QV�`�5=ї����hI0�O*r�^�[f�θ�Ӆ����Ö�M�C���kZw9�m �i��޳N~�A��;:^g��A�{Ef�J{�4;UNXv�4�R>/N*��@;�#uJ��t���i����6�vuS�pT��{N3�-�*2�����1���dĉ�˓pƸNy�Ϭ.�d����0к(va�,Rnu��!����a�#�C웲O���B�h|
0Q�p��~�ay 6I�@v\��VZ#ϫ��vW��p�٪1?&���9/�谡lOx7��+m��~q�")3���}��1��H�*��û����S��q�On��Ӡ�	���~�����( 2�!���b��~mœ��x�S�^UXq]��R:*�r������aq$(��#u�zXL��s���N된'�]�і�1Co,).��qCby��N���G{�Y*�O�)�j�<ϸ����Y�ũz���?M��8��݀,�� �_�edނ��� �E�;����X�V�RL_F��d�~t�ˁՅ��Җ���^w�{*��Rd�B#�	WbˏG�%FJZ����C�(��|j����x����`�x��t�G���'�|$����D�C�[&ķȽ��riaO7F�1nXc;��Oj�#F,Ab�Z���2���=Hm=kM����>(61;6#��j�5�u���킥��y����+tufz�8ͧ�՗�7,����� �����F���J>IаT�5Id�f�g;�l���O)q��Ot`�^����Jb��rk��>K��x7�U��Wbo.����k�����Y	��RM���rI��a[צ4"����
I�o��-~'�7���!>�h��=�\��,�8�G�Kd��Y�]q:�kǜ�Z?r�E�B�ȫ��t��ä��9�����1�\�w�­�_�ܙ�	P]�;rj�/��fw�ZȜ�i`����Zs6D��?�Ζ|��f�~Qd܋���Z�����O�N�B���F˴�,����X���P%��w@���w��7������ �V@%�J�AD����0�r���-�2p-]?����w�$� �bp�D�;.-�J�հ�%�X�.'9w0ɍ�H!k��k)?,t�����؊t��eS���
}�kq�!(��̥������^6��)]K��F	��w�D�F M  G���%�Ғ&���ޖ��q<=�u��|�Ty��Ŏ�ٻi��>��|!�cg�4b� $ߺ+��':j;z����v�+������ciХ��x���h�k�����Tě�Zв]�CYT'H�f_:W��񝯅���$-��fRk��`��re��ޒ�����=�[ �j̖cC,��q���{��II��c�����<޵���Rڤ���:�2�͹���+���붟�3��.�;���}k�P$ɵn�P���s��l��0sn��osH��C��ʃ��Zy��T͒s&j~q�&�z,��`��yLƠ�|$��bL��a^AI�Wa�t�0j���(��o����f������ؑ�!hd��C/i�kEUf�W��N���g��D�8���Y��b&[�� BC�u��=��W����MrF�k����J�,	����!-�S���m�s1�O��wd����Z�*�i��Zz��ۏ�x�+ҙ;�ہ��.��9v���fuwn�q���fE�P��^�0�N�W��@��կU�@�]#x�gP����ڗ�fί}0��,�7F8"%~�*��4�4^pI\4"��0��2���������piI�c��/�g3�v�o��_�#����F	��.�����"���kY�9^����z$�l��e\�axR_0͂7oثc;o����t�S]<�������"_U��p�eb�v@DBz[K��_�n"�P^�3�ì���J��-��ퟆ�g�3�J�KTb��>�p-l&���������%��&����6ٗ�G��c,�6tQ���d��,{����Pc����uo�o¦�Zƺ� ��Ds��3�!K�Tk#����s�������*9�g8�{s��׆|.����GK�Fq�Fr�H���8L3���̈́�y�M�w�ܼ"0���Ҙ���c-z��$�iK�̺kS
�7��l7 ����Էzv�|J42l���'�5�W�{t#�8j���9Xݬ7��0�m�!�-EW���)b9#𫖍\N�
gb�1��^��ri
�2@ڌk�a=b�M*��7Q=���%���?�)N���0aOу���6����<3ҧ� u�x�?������Z;����\(`�(��Pz]��;�?�K�2AWV.}6�;�a�>\�9�d<Sx��4��><��s�M��۹�d�֗�.XR�@:�y�љn��U8+F��!�m��|�ϵ�ܾ���*m^Ίǧ�-W�}© N�S��l:�������F>�:.�4��$�Y��#W��7Kx˃z$��j�.�Km�4���u��u�n�Z-f����2�~����x-�"{9�tQ�p���D#��^@?�ݸqI1{oP8�E��n&����l������;Q�9��v\i���G܃�/J�9�ձ�H������z�����a�g��Ȫ��,He���@Y�j���2p���	}:���w�qdL�Y��R7;�̀8�K�'�s/�L��,Cu�c���e�R�W�6zS���QB��<�f�NuB��X��Axi�iQ�e_FH��]���8��\ �Cƿn�ٖ��@����e�:}�|g��E�Dr�K֏����(A��&��Љ��Cv;��r��d��k�����c�#�bu]2+'!A&�+�rF�@9�!��1��KԱ�?��n#����xYR���I˹�W���"|�$��A��0^`<�;�����>���%�y?R�����4�f1k|��s�-��%�(��-%%��Ή��`�r\���[����\�pe"ZHy�Ƙ�l��3�A�i��t��|�\�:���,�=	�B � b�=��L����i1�5�rȥ�߭��_}W��&xoғ�oD6��и�+`~U'R�y�Z0�K&9�&}�6��Gw����[��KfKt�/��c���C��֚J��*�p+kt>��C#O'�����$�x�$ʪY�]�nϏ�w �Aѵ���
t����]�l�o�/MI���{�jyO���e�4J�,h�}����'4���~ND\����b��QԚP� &Җ9���'�K~"z�V�Aܕ�2w6��3�d=T�*M:�5틢�e{	�[�A�@��rQ�B�&Ec��k������2���ƾ%�3E�L��I�,��0�Dґ �� ����IL-e8�T����E�@Sӧ��p3�[��I	��+8;WS�ǟ���J7U�C�q0- N����ݤ␴�Sg;�!L�	���ШU-n���.{�'G�����x�Mjz�q
��<�Ii�=�s���*9:!3���~U��̇� ��)Q�P<M}����^*��/f���y���Wv��6ՙ�J�1T��[C'/#���t�5LCpO,��m�3i�gv�arEy�eê�'����@� GF��m�oQ4	����&�3�!�d%px�0�8H�e6�}c5mI��bd�$��>
�U)j��	�������@����K�l4��9�kaa����E��3S>��
|�{��tE��O-<�y��1͆��&L��$)3����C Ba~F��ؔ��X�x�(�<_�=/ޥq٭���(h�$C�R����[w}Z�o�"�9���zvTnZ>.��t����na� X�v�M%��U�־��:+#�	�v���Ϊ�$v�ǜ�o&
��$��}�����2�㍖'�:!eA�ê�L�%�r9����{��Q��;|��^�~�_��Э��Љ���ъz�4k���6���z�2'hp=
�`C4�
xԔA ������M��������*��C/�B)����kl�.�Q��FWS�6PC���y;NҰ�i��L��"b�����V,�Vh"?S�m�(���X��k:�1�ҖQm����P��|H���m�t��[��%���f/j�3��V�m�~�N˽�����BG�MZ�&;�r׼��!�ѰF[��j��P��-g��0�5���q�a� v�h"�T��B/ճ�|�+!�Nl	�;���� !L��sK�*8tB��Mʦ�������ʳf*.���9�@R����f�	(��x�J�;��DkX�89��%˄3�dd�TM�JB��]���W&`ۉCt�w�r����*�� �4u ����cL/2	����:��1R�5��6�s�.�܈Bϴ�q(��+@�p������YڒP}��׼,.)����MQ�e���ϸ��2|��	�:��Z$A7.^"����J$�6�:�]���$qQ��[4� �����_ũk�4����[��i�UB�B��9���Wv=$�o� �k����\� �/��s�h).�8J�f0���~J���.)q�����8��
��nY�^�C!QL]k����J���ݠ-Ӡ����r;¢ n�^�h����5%JKӽșO����3T.��?��	I9J�"+��؎�����߈f�B�y<���?~�cX�mp��ǀ�B����i�J��j�0|U&����t������7�>��s���-Qb��X;���r�5Vε�"<�� ���+�
%���}K�{eB~�0U�P�!���k����YR�U�c�xX�,��}�y0��ߐ}ߢ��r(�`�~k`�yr�<�*�F��C��Uܯwq�ۇ0�|�4Y��Co�yd�I9�"~Sү�;LU���X�"fu���D֫F�u�^^���e㘼��k��W�U�P�¼ț��EX�0$������ kDO����?���y�찀����g=�C��=tD��TK�5S��ڝ�ý	����
���,	d�3��^� .<V#����%�RU�Z§�e�G#���e�H���y���<�fƲ	�!2H�}�1�����A�AF: �yfg�s �����U�xf�kG?�+�})�܎A����J�Y$��B��e��W�9*�/g.��QR�����T����j���[�UvY���7���7�d�Qo�A�mcO�L�\���G��y5zc
��0-�U\��'������<�"v�w��GU�P6���}������V�T�d9B2�n�+T|o4�~�owC��L�ֻ����X8������rbo�"긣��)��Ӣ�mo�iG'����}z����:�r�X�k�M�.��Uc���
����ʤ�1�-^/#���0J�07Zg��D�ُ{����{��K�Xᣑ� �X8�=n׫�e��Z��N�� ��Z��g��_�;qB�7�L%�s\��	�N	���2��mY�#��O�ܟ��b�'!��.���V���$ݎ �����.����{ȁJW_��$����)6���� 00.���y={��()���G��s�h� ��Vо�q�ONV���`�!2�3<�\�bf�0�)�TH��ԟ���SCu��H��9��T���I^���J:&B�,����K6v������D�V����O+�����DMH7�Y4&B�:zӋj]@҆�9��R8m�j	|܁ ļ�,�ӑUt_8qbW0 e�m�<�9��P�=�[�d걺��3zv{�p��aV2��=� �����~�B���ՙzZ��[�c��b6��'Q��N�� :��.�D��B�����B�a�b�c�W��Ű�[��m ?�U���"7� r�Fh�#u�<�/��G����稸�A�,��|R�~�)"k��X�~h����Qf���@�+�s"g8&�EBʴ@F'=a�S��w�ق�Ok
�9�������^�Bv96`�(i�� �*� ����B�7���[����{yrnN�2(���A�s�j�%���DO����֣C�LC�	3���,L���*l��X�2+�u1�A�y��a�M�%�s�!ϱt�y�9��㱧t��H=*�k�������m,��Nn�іvs�?�|�妉�K�u��Db���"���K�jߡwL��u�������Ň1@}��C��R�((!/��7���(�w����Z��3�j/��8���s�'��}؊KN7��F �K4�{jCs�Ɉ$��R19! s1���Wʻ	RcJ����|7ԥ-��oM3M��m\��e.N%������S�8����A�B�gKˈ2? ��1R � d�X�Z^��/�FF!:�p"�ή��GH,�$sW�B��u�n�y�D��5wk�:�n#�o
v&���3��[٪xZ̴��@�I�"�e��}���C�O��[�sS�v��/���I�:�X�]K�[G"�U�<�b�'q�hu�$�R̈́a��]�q0�
#�߬i`8��`���k�F�uV�T>y/C�� ���q�j��(6( �a�m{��X_��B��k{T�j��(!R`ߖz�%"O
���n}�㞣%�PTt���hnK�"��*�γy�/�&BQ�����/S�;��i��l΄�&+ �,E����l�.��x�v�~��f�lԞb���G��lc2L	��c[�5��3^�nC�ʿf�d����ze�\m8n�\���p�:�C��C��~Ve���ܵ����K�ހ�P�|����s�W�x4��E�Ko�3��JJ�a�YzU���o0�-2�p���k��(#GN_}�=S����{��XU��T*�1C'�J N��g�'�K������ׅ�W8G!�Ƭ�e+��u�`�uIf5���ZlU@~p��u�W}rU{��a�;�A����&�
��0�?����5�1�!8�k��C>�@�nm�Y��f�K�����ͼ��7�:!�dXh�o��10[�;����^�"*�+M=�kt���כY������������2�o�� �E0X\�x���;Ա] S�
T��A��Dw���+'U?�ș}YM�����a^l'Ə�t$��Z���rN��7�a$�{�{�٦��������}�>�o�*�5g���EY���oz:�+������2�1��G�a�i
���h�{7�0��(7�ۤ˪�zZ�t���.?�=]B0�(q)No�Eh�*�7��(�������ZLI���f�置"�Jڒ<{�& �U�"WJ� t�T��P`�?�/�~�5��0��gLH��8��"�nw�������{�#/�������q|�׵1L�砚��x.��H�ݾ#�UcN,�p�T�5I��=���R-il³��	/Ǽ�E�?�I������y�64F�lxj�g���iDY+��X�ԖH��R�Հ�Nl`�h�q2�!�����zUk���.j΁������8�q�:O�J�<�`t�E�h1O�����|��̖���ف�9�!����rRՃ����j@MÒbO�Rʰ��@$2C���*`����h��,6:ݍr�Cť���6d����E��0Z����3����w�@؄6J�埳˂ŗ�:�%U'��4"\��2Y�&t34��<�h}�$�{Wc��ֵ����'�!K�dksu�uj����]\i�c�ɒ��֫i�ں՛6��+(UMvLb��9�fe��wO�1�kت1̱90vO�_ݹ�C`��{�I���xqy��rA�3�1K �K��N�%tx�x:D��Ϸa�n�>4��i��B^@�`B��x�LсD>�w�;�6Z���;Ŷ����/>��Q6Q��.�8����n�����4<���3�t�׭��d�ŕi �L6���5�2��+�W�K�<pH�++��V	����\u��9�^s!Q��_��-Nvǜ�y\Dg+���4��T�l�{U�%�����	�ί�a�G��7V�`V���0P9X�n6JH%��r�=z����ի}�WuF_s��E=�^�5����XBuX���Yl����#�7�
�V�f�dmg���o�-T �o��M�37�+�����������q������_��f�K(✯��� zp��j,h�w��w���DM{�7�wo��wf���5á��k�bQ50sS��x�2���ՉR�[G���{�Ý��
̦���\��R[��`�$��T&�C���B�e�qb��	6�����Qjay�x%��F2E��~q�	�#�t>��9zFR�MN3q$����BՈ�L��HG��j��LŻ^Zo�GL��8[�L ����1h+BiY����z��E��%d�7f������z��;�����<P��!�)=��σ91�ቦ��7���N�J�M�'�Ps���0���xrjY�#>���!v/�-Jq���;u��-�X��7�x�o�z<H! 3�Rp�_����48+�����*�'�j�l��M�ص�P.2�'�5j�n]�_�5�W���B=L�s&]�(�壽�n�󡲪K3z6 ���'m�,@�%�eĤ�dp��a�Vq���@ #�f����+�9�\��n0��iy�rm:�j�`��9�:�INr[֭���BJ��?�ե3�N�l�U�f�`�#������z5�f�ݷ��!
�]]�]�+�V9����3Ip��#
DhZ�qh�VZR�`��8s=�pkT�Ȫૈ}$�d+��*+	(�w���r�y��F��&q$U�����F�1�j�w�Lj
�I����./��3�c����"��f���Rϓo6�>���"	����0aݱ�0V�.�%��ӣ���=VH��gv��,?;|0�K���{[�uI9E����ڭ��H����@��'�G�ÃI��R
�q�
��y&�oP;)�.D��e�{�bx*��[�^���Y�������%�m�,��V�qF��x�`�]ZW�
s���t�,�Ƀ�M�Z��U����D2}��v�����Q��i9�]�ki	��ܒ;�ʇ�	�Etz�U��*������"���"I�7����1����m����a2.5q�ܵZIV:��,�L�=N�%0�%jm�� �4�k;l�)/��-R�Quҕr����fB�#��k�E��}΂�N�*�sd��*����lo��T��$�ֽ,&�_�����e�$�
�@���B������Cq��kъ����F���'�w���d��䛊���Vw�ʶg�S+	�t�o�e�)eV
��(���e ������m橓�l^�V�sM�֦-��J������x�1	R���D�4s�#f@��D4��$o�)�d��Y��D�������=c���C��/���.���?����9��s�s��(�B6���:~�%ZsA�'�<M<wRZ�OW�HO`��7�N�p#�5MW?Q�^�lj��PН�CĴӣ�$t����Ŧ12gC2�^	 �����`���OiB�l��UR�A�,�%:r`t�~��eDMz�cz1�I�*��$}�G	1������+-�éN����W�g�Bp��/&����"�?~���u��P�iy�6"�TGBŦ�-cӕ�vE��W�E�U�8V
Ҡ������IS�k�a����Hf�;vpL��?�*3�����}���w�6C�'X0�B+�g��V��'ShWoƧ�⸎zI�cDöwu�KZN��hn(�v�P{O�-k�+�%�� �]��a�vk�ئ��s;(\A�6l��jl��2�>���L�5�	�n�A���L��MT_��;p.W(*c���
8
q�����N`�TTܾ��Ój׫P��a葉��)��	��*����y�͋0����T�HE5i�*��Ê6
�W�p�%W��[Y������P�n�&��R�mwmC���51��am�q$�����y<��E�K��zV��ٻ�Qޔ��"�SC����pѻZHܟ5�����$D��$��͚ko��F��'+��m(�Õ���魧JY ��&X��,҂Ť��E�"�7*�c�V�ߣװ��c>���5������u+X���>�y���I��\�7��K�)bƏ����C�LT���Z���}ed�F��h��[����L�k�\�����= #�9
]����R$��d�5q5���$�[rs�1�Д���Q(k��\���dX? �����^�%���Ϯ���f�}�K����'���������0-� �A��<Mԫ��i�����|k0Q�c�e"97�k!N3¦w�7ϭ~�.�-�n�RQ>����iY��ѡ���S-�(��q2v�F�l��*ۘ�I�ȧ�#�C��n���>D�핵
L�U�jW�q�Z�MD���5v���1��J�#�櫈��%�TW��0<Kחw:M�ͽ��u��zmy4�({����
�z�f�2���킟�o��X}is��� /��隢**��DQ+ �^ �R���0��ƃ�lc����H�:���4�+u9�s_����\�z{&v�oU�{I��b�x���d�>���d�,��4ܗ����ݿ�\*��J���9���l����}�×�yL�V�Ro@�z�>�5���	|����r�1�QF�|�02���4�rJX#��p@I��l�F���x|a@��h�Uk�.Pd��H.�Q���cƏ��M�#�\ceP$�ARC����x�@tsk~U^���l�Ǘ 1|*�śj��-��l��(C��s d�;*�}�$pEwf��.t�ލ�|��.Dʑj�w2�) ��L\��I�� ������?u9N_w����5�MAF�3�8�'y�B���?��G�~��?��:Rc��>!�E��zRK�{���W���vl��=����a��72H?�{���4�c eTJ�颃p��榳�g��͆�kr����OUC��W��}�e�oA�N^jMo���lSh�X)�kr�џVom�������ܡ�����u�_#bY
���:lƧ+���Q���I�D��pq��xXi�1�`*ͻS�+��'Ѝq�e���ӻ�U,r���dy>��b�o�<���vfPDw:�A>�:�k�u�e�%Hy*peI�X�Z���i���,�3H�#�_9��-��U�0�l���F���;Va�i�m��.��J�Ht"�n<�-�[�S���o�
�a�w���i�@Y`���,�*��(�w�u�S�è���x�\���H���wǲb�'�:��
�K�&�"ko��H>*��{��-�p4=�J��N��^T�<��S�
�K��m���]ÐY�V�Hw�����,��$T���#��bi[�mB���/��7���
A�`<�ŕ�U�t�v1��s:�t-7d�U�)��mu����+{8 w#�_���s���V2l��#��Y��6��	����J�Ծ�aL=����!�п�&�ܢ�)s���6����T�W� ~>.��zp3��cb���X�#RM���<�}G�o|a��؏��c�@J�s\9�ͥ�*�3��ҰZ�����iBGڹS�O����M�\jd�c���03a�(^H?{3|W��j"��D�,F�(�f
�7�<��*&A������ rn>� aj1VG�=:f=�3��r.�^O�):5���lv[j�}/+�>Q I�V��I�@���|�3҂\,S�B�z���	���f�z�U՝VcL&OX4�!�FV�88B)N�sZ�"&�����+��~�x�ȡ���(����!����tϦ��fjP#(�Wrp��9�'WX��<�;�|�E�b�/u����H;$���`��Cs�>�
(_�}P�!�����A�9(t�Z��*T�|�ͽ�+���~�~Ń��
������C�������<I�Z��:[�x�^a�YB?�m�ʷ\���Z[iMP��^�rd�ۉ�o���<���.D�_��6l����vÃh�Fj��=��s>{s�L���Ʒ��I��T��,^�4~��~ �=��+�F��Y���(\aG�g���燭��[&�OIꡜ �$�n�6��b��N����*�ߌ��E�SwFEH<v�ր{W�����\���+t�+�������+OE�\e��4�vyJ/FQ�$&�m#{JO���A�=#�z��fsZl�k㡧�`"E|_ ���5p������qж��HPK��4ٷK`��J�x��Y�g��se�k�1���Ƨ2�t��Ǽ����J6�3?W�tm|@�����<����T�iZ��3�=�J��q����]ƃ��M4���t�=�K[�۷��y2��b�T���f�����|hP�
]{:���Gu���j�rW���MN%��|�l�X~���K��S%�7|7ȣ>V*�!���Ȧ���&�4�A5�
����.�*���.�r]�k�!:�Jε%�<ҹlp��"�<rh��R��;�7D��K���e�j�>�xWmy���6�w��F�&���IK۰S��U.��"�������Q���΁#.��4��I�>80f��PQ%���ƹ�u�Z-+����d�� ����8!�A�E�����[����<���S��A2�ډC���� ���J�) m_�aq�?��Q�XXk^��K�#0��D�����o�.A7l0��A�-H�3o��}��Z
�D����b��
���E��#-�ë��Z���DRiͻ5��5]ϱzn��ì�5`O%�����
Kɤ7Ȃ��q�P풆y)h��ϯ�(������,$j�H{+��^K`L��6]^@�SV"B�hL�S��+��=!�I��P����M��3�����b��8Ӎ�8�>���!��׶���Dq���J$$�j\M/׏�˟G
Q��U��_�^)/���;��4�"ky�㵥�����FK��"N�X���]Swr�d�`���U_̔(��xؒU8�<��[K&y�36�*]+�����%�i&XR7�&m��[c�X����&8�J���l]��>;��R!�z�[Z�IBa@c�,�^_�F%�NxZ���� 7�R���f�+.����򃣿��¹	�v	:c#&D��@�Wݧ]/^]��V k��\�]���[:O�;�hwv����P�k�<�EQ�X�Ij�m?�̃�L�Md@��?��~\�\��D*!]h��M�8��8?ìө3.0v���l-���+�¼b���VBa�;<�o��܀�h�ܡ��~��N�><j������)<(� T���^��}%m�_�ݟ�s��K���ѻٖ�#�ڸsM�ds��ެ��7�hF_K�3�
�lx�Ϫ���q��"�����?��ǝ���ȝ��d��I��x��tC�[U���*���;"a�� ��G	���H�d(|�jI͌������q,���j|��2�X#�I/5xChX�mZ�hD�5]�󻆮՘������;B�q[a\�������S6���,Y��p@�)/�pM=5��G�S�'�0�x��h�L���c%w�Cv���S�4�1��ԀV�P*w��o�E�h�GB�Z���D���)U��fF@]2�b# ��U�뾕�C�wY�ߕ D�zZ8ڦ��mj��	�����"s�F��?�L����@��S��Oh�П�-p��Dźj�RBӪ}�!���ѿ��(�XP����}�'�dx/��dIM�5�zo��S#��i<���u�2*��)@KY�褩����xl\���8����hK��Ǹ��4� �- w��ˆo^֚�?��M&l�����ha���T��&���MD\BE�5TS���[���隽�~F��e�"�����7yq+��I0I��	����ړ�������j�L��+��V��%ݔ[�`��0��{�!�3ErЍ9�^�!�h�VBJ���f���D]q:4�N���Y?a�$��ܰ����N�(ȡ;����FϚ�E��D ��2)T��}���.%�A#��� %������n�")��!�<�QRg�}�m��(%����Fp��\�.g��j��&��W��Ͽ����J'y�K�0/�V�v����[��1�#�*�aL�(��֎Q&��V06��X9���-���T��ex�p��ݘa�@����Q֊r��)>��t����
�'�Ե;�`�&Fl �Q�F��OΝ�z}��l4��p�B�K�YX�	'�v��u��j��=ӓƀ�&��t�re��<&�����Gʚ�nZ���0�{gk�	���=s4^�y_��?)��B�$�;�V�rYBY�O���\0���Ș��
S�@���H�ֲ֪��
E�G�V�t���duϺ�2��#����=����-�\zd�Ǻ鏺�����&����h�F��Ix7:e��	�~��+jG9�xB�'��X��1�[`A@v�.���d�7oc> �`QP�i��{ �7y(������)d=#�دi�3Ծ�U�n�����c@��I���$���&�h���<��n໱n��O}ʺ��v���)�����<	p>s>äm��ݩ��)���Ɍ\On H�v~}����0���	x��ť�g���,c�)!�mtNm��4���9F8�B z���GL���rm|hQ� ���+_���H��˳i���vZ�����c���x����Mh�_�7|�SS��sh�0?~ь%\qk%���F�b�'<��?%������,��=���v�3^��lȭ�O����w獁��B*���cI��#�lʙs��ґ��0 ���f/�������cH9�"KoY�XP��`Ũ�~�i>Rece�;�nL�O�[E���5�[�q��t���xyn�),�@�ja]�K�%��MV�!�J�#���Fo&N�q�ߣHu�%�M h�i����������z���D�X�(�4��k�����>Ap�R���*���9�r֋s*eT�U��ſ�_���4��G�mƺ�R)��ĭ����'~��A�pA*̢��:H4�$[/�׷�f]��2i/��#B�(�.�{4�ं��Ro�f�&�ߙ����d]��~�c�Z���>έ�E�#�z�g��d��i�^��T
����e�ŕ%�%m�Մ,��I5�$�7~o�a:�|�,��_Y�F ��Wa�8���\��Y��|؆��8�_r���Q�[t��Ca!���d�2(���|�6IѤI �Nu�(��s�o{q.L���%��*ۿ]'�?�,�EPy�n# ��-�rB?�+1 ���e�@�	9�Ӌx���Ԝ����n�L{����u�%R`{Tfm�N������u��z^�=��/��ǡ�B�2�S��}�k�7s��ƽ�H�rh$X�rqv�c<hJT��AA�p;9��wRM��p��쨒%�}]*O��� ��HPqP="���W1i�<q?���]�i�!�]@�v443��8�U�tȜ*�4�Q]��e�@�S��K��O�oF�+Q�5�Q��A5�8^�?�(�	�>���O]1��ݿ�;|HR�lt�䔪?������KJ��妋�;��B�4IO��u���zu��[�1��.�Q����n���zI')ĜA=<�e�3��d��*_��@O��R��-�7�f�
��EM�Ggl��!��~���j���"jL���m������R�J��_a���z������tU�|�9�T�p�%�e�U�p��n�j��4uh����ǁ~���s�p�}J�"���=1�x�.��:�.I��G�ߚO5ܫ!*z��31�RR�2Y��K�RJs������q�0�ux*��K�Z1�������{�;��
F	�c=��:��|���0l�L�R�冯����iC2��7�T�^���V��2�E�I�&I��$9E�P���]�~�O��p=mg���'���,@�'�¥��8U�>K�$5鞣o�%�"�Zv�ld��R0ݵW�7�{:BN�����7ہe(}�ڙ���ErH���(�i^��
LBH�h�V��v��˱O��N0A�Ϸ��2:Ө9C��x��VpN���Y�h�w�����?)��V<�����^|�>k3�{.�.�CJ��{�:O�v�փ<��zS���nk'����::I*�`�}$����d���=�5�x�O7��6�{��+ڬ*�U&F�J���[�m�v �?�f=V�(V�gl,P����B�b�����m��($hR{���qD���~��&.�-_�.F-�.C��&u#�!����޻����4L�)N9z��6��p�?���x����q����O���θ|px��S�ɿ#��]\�I; �Xod�@S}�1Q�kү�L�k����Պ�ci�S�J���e{�X�NH,��$��
�ۢr��Ku��� Z�Т�A�0����-�Q�v;�~9TK���K�N�g�T<7ؼ:�m� �������?W~B�G7䝹��<����0�c!��VvBU�[�6Aa��Pq`E0h�6F�BA*�F���l�����1�u_���!����=�.��]1��B�y�Z�N�B�N$�چ�D/$P6x���<���j�L����Q:�=�}Q��� ��&����Yg�E`"�H$�?.�'_�I铯��O��H��Qj�$EG�*^Z"��	t���ٰ���0�ineF��g�gŮ�������m��[�1vȧ����(�7]�S�2�PN�R�e;8�1o�6�B�(@(�6��y
��3�3���3�~XKH����*�C�ys�e?����mD;��sT�%�`���T�Y�J��TX�Y�7z!U�m�ב���v�����Ooc���%�e���X�M��V(�Ȩ����j`V�cM8��4A�P��� TSW�P���)�u�d#?����v��M�D0�"�T��3B��V�v���k�1��+��Bw�Z�����C���꣒�n+>�#~�����'"���$=�};[���:B~��F��SVs�Fs�}k�
)���8�Y��1��E{X���_��q��}���[D��s?YB ��=\.6����W\ѱ��C5��8%H¸D���P��sF�x���}�C��y��F���4uA��-��,ʭ���+�4�$�H���m�jf���y=��_#���hmwѠ8��]1�n���z`�b�����'�����r������ u�ſ��v:��Y�	x�'�c�{zv	�iO:R[ei���E]-� �q���ߓJ���7��	�҅���lttԹ\�K�J��v��t׫垖�&��;�^OV46wT. ���/a`�}^�9�"���ߩ�DE�g�2�aر�����2>�H�y�H^��_� �$Ac�`�VzLSu
��:n��X櫞bm��	������F�ï�`��1;��؟��a��p��Hh�7P1�NH�u0����˾�TP�,�"m*���j�	��ɣl��셺<fF���]~.�C�H3ҩ�op�=�;��҄�����(�����z=fV�H���WũoHa�z4G�P��,T�ǶXp=�̓w$�l�VAEs���Z�ꍄ���oE�࿴�<�MR fET
R%�
���J�;t��b�D�?�F��簱$'ԀK�U]�a�����%zuXy���d��i?�z+4�(��Cy �p�i`��<��:��T9+��+V�H��O��#�`���	�ɌF��C%Jc���R�a~�~UQ��6p~R�WE��9נ��<1�VE/�u_c-�_ǳ�*�AyI�
R�UH���u�oJ�Fz=?�����$�]��Z�����a,!]���p�D�U���zh֕�"</��//�,.,#n�#�$��R)�Q;�,�#�3!S����u˅�frpo�ɞ6��r9����]MI"E�?zv��M�>C(�����'��SB��	o~����of���:"'h�����p/As��=�ݔ�8[孃����F��Pz��;��1)�A�ſ{��kT��:ED�(Q�����If���rJ�ɕ�[
������dy.tH|p*#
6﹙��/I#�{�f��d$�������O�oޝ.L	����myt)�Q� �������Aը7���y��������h+eX�{X`�8*�ۆ��}��_�R�un�]��˰ש #"�˿H�rبv�H��T���wZ�C��L]a��p.Ĵ&���>Fq��{ƀ}��Tp��w͟��V��jEg�i�%���f�P 1^��|�L����M;��1ЉZ�h���N�����[�J���Q����g��3!S�&Y����|��!0;-`��޲v23����]�W1�%��H���Uci�JX�p�z1Fc?|]�t�@��Id�&WR�t��g��Q�|I�%�*,Ƚ'U빝[�'���*�l�1:j�(d.2�|���Y@��n�"{�tK��g��u��6�U�&�[.\a��w��1�g�nJO<��<*�v�R%J��
�^�x�����H+!�^<0+���b}x��l��,qKD
7W�UD�/�KF��H�F��#���]=�Q	rX�\s 6���lF�W,��¢�"LP�)T�`��F�e`�冝��#��>V�FJkhH�[t �^?V���~����J;�G#�7��S�����7��n}�R�č�.�8%" �tM
�<��Y��'p?S�=�����^�X$�;�L����w����Pb�vRR8���4�r0���;�퓣�Y>e�t�����%s	P�w�������Y�?T����Rt4�(�q�U��Y�i1((��F������F	�t�p���u۶q�,��J����+b�hs�`9נ���z~ͨ��H�eW��d:I�"�!�ڝ̖|4ww!o�--@�C��k�$$ȶ
'V�$:�&Ś����+�&��t��K�V<� j��)�X����j(L�Aek����#o�^(|��Q8�Lq.�'��i�b����t��Ju��Կji��
ib���'�*6�߭� �$���P�`��i#�H��ʚ�s�	I��W��\��V�:
U�pA��|��.���f�|���� t���x]��qvXܵm{6L��Û�EHb�W5���bۋ��֙%�a�`EU��"=��+F��y�}Ո�P�9��P������RY�݀���#���'��N��F�v��8��ks�nh|DP�y<�ӡ�V�3�J1��;�� �@����1�P�A�>d3��߷�mtq#�l��}6�zV*�W�0�[�2�7�D�ǌ��

�>�/ K>pA`G�S9�B0Z��e�k�|���&��K���U��#���X�K1bˑWՁ���ϛĬx���"K�ux��gs=�,�8C�O9%�͟��vs>�2CLP���́���k+k�W�o����x�WL�_��5�W�������j=����
Ҕ���vs��ᑗ�ko��B��=Y]u�@��@q-��/-����&�jO��T��9{���2O��5K}?�d��+P�%;�ûwZtCͰhmlf����a��@�Տ5���x P!���1�����������*H6�rB.�������U�<1�����%::$�+Jw?ڹ���`��w\����!Г���C�*$w��A��9�#��tT���6q�����G���ʨ>�.P.a@���a/�>�<��L�;�� �+�`���A�y%,:���|��	�6g���@h�R�׬�I���+�����[_�����'ݩE�)�k��dO?�裪BZ�#�e����p޲F�`Iih�O��=M�T��% �cc_1V�|bdf�F��fQ��b��gh��`|'�^4xY}�+x凫����3�2�ݧ#���jd���Y��8M�Y��U3���,ɥ<#�,����E��\�X�o�W�E�|����M�/�z���?Z�e�#g]I�y��� ߺ�39r���LQT)���) 2��2~Ɣ8LL"�Jl��͊SB���ʸ'b�9'`y{Q�؄�w�f.ҹLG�&�o$��x�p��F�P���Wn��'��T2\�:/5#71(Ǵq��>��^+v�p*��>7����m�|`6x�cw�	}����mbfO���٘�&����'�Ml� e�Z3�����[�[���ۘ�z��q�f��ڹ&D�d���YiL��إu�<�h�w*[Ĳu�.!� �ǈ~�=^�KQ���d?&�+�L)�v*D���u��[�|���}Y6
e�4˩���|j�ay�2Fǭ> ���cܵ�5�\��.���0���Mv��dv�(%��p�~/���>����uM�9��q��|E/�ew�P�f �h6�Z�Lrǚ�.�����RD�[�L4@43dY]�3��/����Q��v}^x�N������~�?	�Q��;� ���up&��rJIX�2}��㐰���n0��fe-�I��u#d��І���鉬�Lub9�񅛡�c+Me�����U��wMw9�su*�\�� ��7�z�
&�����3��t��+,XX���d�b��R%��X���R�
m2ӫx�J8��K�󯪈�zk�y��J�W�X��y�C�%�d	�Ѷ�Rj�<HO�R�>DSmP�{�Q �i��o�v��7�u.�u�A��<�n�x�r���b~�V��b=<x�K����y���iH�"g̾*Csl�6Cd1�H�?�Z.�@A��1-M�H���䈘xyF�`<�aSv�e����x0�����%��2s4zXն�:Q��_�d�3���K�]X�d�Ex�EB϶$^Dm�gcg���&��Vع=��gxh� 3U=N�.;c� [�b���'-G�wG\�5�9���Gk�e2P��j*��W��|�FĮIn{�W*3�;�YĲ���KYсK�,�θ5<h�*��h|��Ʋ�/�b�/Km�O쭤y�i��>��r�S���Ǣ��;���77��кwO����ߒ�z@�87���o���!8�����/�ʀm�T�a��;�fur�Y��E#�l��-i��������Gt�ʂJ������n��xd$Ο��ǹ�	/�ͷy�� u��%�Woz�V�-\�S����.�>�M���.���5X�D��R��QT�zUF�T��!b���s�9^k{T��	�oF6���e .��8+�>4ۯ䙛��S�Ata7�){��l�a'$ۇ���E;�%_G�[��K��`q�<J��*�H_�J��x�<u/6*T���~��s!���<�!S"H�u��^V��-�X��AxS��8R�����5���7��6�(\ERۄ^=���}�{W��4�?su �&�F�w�D/]#�@F����-�3G{���&��)��#��K z�dvh���>g�r����V,�0�l�!�&=k�O܄����bw�<�]��ڣ���X0¶����"�p�6Y|�V�HK��*]���u��L)o ��xP��Ua�le�f*�](���($)�lp7%�`{G�C��+@��%���n�/2km?9�qy�5�Jl-�^+�#+�!<ܼ�X�{%�\���%_,�5zv��yv�QR�ȓIz�-j���O:=Y�5�>[@J�&��5�����d���y�]�ᤵ�9U֤W'�>���$��u�k_��$^�h�?hU�ΔY��7\���M�)%�a��Wa]�x�������5�"@��;B�D����A��g���c�@Gء�a� g�#�R�.?L|�� �M�����ѶJ�]�	6'� o&m	���uv�t��z$A����0�h�S�PR5i�O5ؾe-��}â�=S8����P'sy��(uRkM�!L_�
�xlm��/��
tD��M��t�<sE$Y'��u[�����fK�V��۽Э��fi��A�������j�����Z�y6�Qq�B��W"�	�*B�����ζ���i;0g�o�[�z�{�z��2z�Tx)�@��'샊�ʹh��V����!��v+v����æc8���D7�~{Ym���\d�g'R\D0�����tP��{L��JZ(� ����ٌ��[f�k�o;����n�K�T.d��h�Ɏ��j�	���Id0W���fG?�J�<HRc��\�3 }��8j\�MY���,d��8��1�/6��G|�hk���JA�$�v�f^���[UQ0��U�W)Km�}uK���uzs'�{�*�b˒p�f�V�5a��%W�%�����F��X]����(s�rn�4��kY�^�W�����s}0�@-���'hZ6>�_y(�He^~��R��`��--�����<�Ճ�ۏL���0��jL:׷}�{��[:dε�ǧ(C��.�թ���V��J���ՙ7��U�K��=0�֦%�g��� ^���j��
�x?�V�"��/��&*X�����b�jW�^�!��6e��������Z  �O��|�ӓ�m%$��zێ[A"�@������\�>ť�U"��-��!��=%a�Dv�؏Y�Y�Q�
����������bYQ@`�7��-�诰�c�?lS#�z��*S��H����>���2D"[��9l��8�\~~�{#m%5'�#���&bi�_��C9���9͇�ma��y�be9����z��8��8�@?O�{�O�e��N����S�h���8xf�]
�z�����56��'߹b�e�j���Ά���P��
6���N�L�}�
O����o��i����K,H�A�C3��p�a�g��>0��}M|<o���@��[@��K�tG���.W�st�ӕz�tݐ=�Q�%a;�q�h`+2>��o`���Խ����tP��D���,��Ut�GGR��t����� 0�k1�t�g C�[\�i��v�j�DIs�:&c���f�@���������2�?\]��&�w�@X�C��'���W��	��8+A�0>%��%��t�A^ݡ+�8��0:�f0T[�N:xޔ�{A����?uSY^��ʚq�W4��tY\��}c?k�d�}d%c�lDv���2>
��dFp @V���KiE�*yD$�I�
�p��G'M���MGRs-Qw�<�]��՘w��m���??���Z�<��h�7ӻ��v�ԈM� �)����zsR*����>�$%$�� �y��ͨo�[�`������lմI��r����{�����H�-���)��nm��`�^���}D��mJ,�i�Ś��*@�ɡ�%h�!�B�(,��B�,� �ܯ�5ɺ�J�����X3Wl�M<"����:4qmM���=x���;��:���8�����J�o�?�9��]��_���1ul��:�J2� $N.�?Td�-E�.7a�-�I�D�J՗7�.����I���3���=Z��8��i�K��"�]�t��������,pI𹮉�3�N
����}A9.�'VZv3�/I2�x�b]�j3��}E����i��E,xo޹*�H�7w��{d�G�ߧi�=.6�AM�T�E���OA$}��N�W
w(���],y�s"ܛŅ�0㥼�\��b�ᯪ�1�i�bw�,z�L_��V��W��w[u���6�d�xd�q���RN���0��9��dT�rv1Ȥ|���d�$Ҍ��O�,��9{޷k���ÿw_�+�`6!Y+����M�\U�J�ᶭ������B-t��y�I/캙$�,_446��#�c�S>�E�C��M�����.L�b�P^�S�_Z,Dz>����z0?�-'�EKr��X쥹���ó&S�mK�8Pya(zO��vTvH��h�l�N>�a�g�J�GM"�u�6����
!�����F�۔ ��h��&w0��<�HK�H���&S���!��I0v�ɡ�q������_��\�3x>�g0���U���Ø/!(^�{W�܉�q;�VKO���c�+��5i@��X��i�>�>�U�{C����n��Z�hu򣕱�h��C�D��p�8ƨ�<Q>[�&HV��q.@�˦���
�aI��t��0���'$���P�+��/��^g^���^FY�5�o�����ŬZI��j�՞����,�m;AQ?fn���xw,�C�Ͱz� �r�x�>J������S���ƿ���p�%��NX�%�:5+��ho!Y�v�0����,Tb����/N{&8A��
Y���L�9��]����`5qd
��_};�/��g����S~2���k{'e�q��*��6����(!0xP�=�8���kd�<'{�%��p�5߮������z���x��g�=�����G������{���<I��
�c�=���r��ǹQ�D�96�Љ�D�V�����zv��^bֳ[�Jo��-�Q�}o��>K��h��=�1��䗊���M�y1P)_����f�U�E4��*{i0v�� 2+��Pw\�j�X�W)ɛKR{�_��l�k�A����d�]c�U5�v�-�	!��oC7��?��.��MQ�UFρ�C�E� M���ܣ�\s$����r���Nӯ�>t )�$�v��N��?|X�HfSz��k�
�d�8r����=����ۢw�� ڧ�g�飄/q��^���BL�3���Z%�qЭ̽}K��м9S�7�9*���;aS��<��i�<>S��՚�nn��V���t�p�|�Mz��!a����� ʩ�	iVw�@�4�w�1��@�����3�g�����[�C����}�.�X�̾�9�灎s��"�-��_�p��@�a�ھ����6����
���O�T��8���h�Y�d�P,㲄���ƁĽWɐ`������R_3:�D���`�Y�QX�v`�xs�+��R��:"���r��%�?���]lZ�+���.X�����mL��3jȞ�_��(�洄C���C�јIgy�CNJo�����X�F?/�~�|�1�,P=Ĵ��p�]?���%-fj��cA~vM��>���#�YG�rTu�
�-	����A�����g��s=s@��=J.%�jy�S�g��k��k~|U/��ɧ�T��w~��턎ck�W������<��S+�m�߿~Emꅸg��?+��h��nd���~31%'J��]oR���" ���{�֐��,U�T��Ȍ��Pz�]>#����w`�e���VT�w�4a2*��W���޻��_G����6�$��Sӳ��/��K�5���]d͡�ɗR�(�n7Aے	d���[$�	�Qr``q�yy"��n���Q����"|��GHb�1�'!.2J�
%��/�V5qfj[`�O?����!��·Y��*�����iz</�yu���>��a�+�4�(I��!4���$��0����~�Ū>Z���.d��k�Բ�!
͸ڢ�����|L��m�4Zqx%P�6$E0uyfu�,�e�<�H���N�ۡ��^�Y0!�j5��-���S}�����hr���Q��n׽� Yq�é����H1���W� (DF>��jՍ��ȡ��0<�D��`�I���;E�_b������.�K��h%)qZ���x�ր�YӤ�m����x�̀�Yq�vEJP��
ZR�k��-N��UBz,!���al�XI�y�l���<!~?N���FD���q����ol���o����a*��<����&�mæ]�݊��n/>���,ǋ�H��[@Wq��1��~�ZIihg����YZR>��	Q&��N^�'c'%_��b�@��x��f�T�Bnv(������d#��� ���:��I��P�����+�E?�.x~�ߋ�j��ª�"��*��2���>OP(�:<��id��;i$�8���0�c�1E���D�Yj�<`(I5����%4C4�kLV~�!�`Yr%L�ƞ��'?G�7!$ +�{�z�D��t�aa�z2$���)fO�۰��i7���,��ǃ��TJ��j�nK���5��TC�ͨN.�/͖���H�� @��Q�O�k;2��NnM�+d�;��0/�	�ܣ�ʈ_%8'���I��/:�q��t8���������0�f��P�=�U����6���Q��|�;�I"D��y�Zg���5��6ª�<�鲖ww�M�������7�:k�A�E�n;!#z���y�׻�9E�z¯�?��U�`\ LƂ�GK����'ݡ��b������:-�K�?��������(W�|�7S�8�?����g(l9G-p�`oVi^��������r�d�N�9O�b��f�6J�J���Y��:�F�'�%�^6)A%�`�����U��ko]�u}%�?Q�)ay�|�4i�ć�p(	�k��#��%R�K�$-A,��}i�uYS��"*�ӨVVX�g�"��
�S-�>�+�SP|��Iq����k��1zə�%@����u�n��uU�w�h���Kٷ�b��H�f� o��FՓH՗<Tߥ�����ޟ+���k�[���W'|�zQx�:K�I	Z��_�a�N��F&eC'������O	�����M<vR)UO7R��w�uB �w~�,�)4�lA���e(�)g�T�x!��C�,���ɐ.��_�vtr^5I���Wu�bg�+>��d�V�d�H��QĔ�%Q;�2߉N�w�l���4f�t�ݗ�ݴsY��U�f�-0�V�9[���h#V�?����< fS�0�8�� �R"����vS*��V�5��q����ᔲA$tAn��D�I�T�J!���dW�������6�p�t����R���?g���(�����/�J:�ɹ�X2�������gX�kD��=�؅��-�{�%��8��R��"�q&t�id�#��CV�S�=��M���V�8�}��@=ތ�z���K����-�?�!���$k���h�uJ��3x� ��W�T���T.�
��?�D�we�h�iG��gJ���&�R�	v%5=����?n��'�k=��!�ּْW����a�˥�n��)�<!\����Ӭ��9�7���.jxŦ�����42��Iy9NT90�}x�^;�H7�]�P�qDN��S-��}�D\8{�D�b~��*��^�xT�X-=��n��[�6�y,I%OB_��:�*;�#/�n���
�p��xp�IM��TwɁSx0���6A�yZ��`�\���}v$������ T}&���:8��#���t�����K����bqP/�H������E�f�����nX��&�Jc��������)n�93���ß�6+>q��90!�ݴ���{�%8����,� ��%����8��\(�@�c�.;`!�)����G��2h���Glf��3Ϊ`�� �4��x&��u*V��Դ�\ǭ�Y?�D�ah�1�w��Gv�ʠ�n�q�R5;NuN�w�5�F<�N�R|���7{#���l�Q��޶z�ަ�]~�d�%ˁ|45��ڈ�Z='��I�5s�pi�A�^�-	�^9|K�=T),a��d�4����͉���p�-�!�GV+�T�Pr�~�E��2���[�h;��'<%��<e�Ygj��-���/����8�Ӯ�TJ��7��(�����~�j����C@u7P��N4��M�^��}���õ��?N���)��j�iE�%�C���w��B�2�\伎C��Q��6�}�ᆳT�>�4��u}3��b�����6��?:� �tWU�+�ʢT��czށ���m�g�<�a̾/�,<��p(N,�����R� �%�q ����hˁa�g��m2���L^�4kJ,��k���c�`:�^���B�g/Wt��� �2�T�=`Xv�H�ߗ~[T�j���?��g$�_���5���_ņ&Ѡ`N�s(�s�6w��#	��˙m�i��&��[:��cy]\��7Ur���<��ߋlUƋ�y������>�a��L�- �O�������ky�~�KI���S�T>��uA�ۭUI�4�i�P�����4C��݂�1�˫��M2����Q)جi��x�qOx���Y�(�f��*���Pc�����hĽ��luQ�AY���sc��	��G��^��ﴑ����&A;��SO���s`��ctCWqH����kz(G)k�������I
/��ϊQ�AL��):� �o��h�;݋/v�&��	���9�܂�2I(4��[�;�`�����?0�d��E~~OX��@���5�ٗ���Д$���9ɧEI�ASl������ز��,�i{ڮW~�EPk�.>;��u+Bi��"�-���.B�ф@z��+�v�w�<ȁ\a�r֤_5��9k�_f��oN����������͟� �q����0J�$g��Cf��cZ�x}L�t�H;0n;���A��]����bun��a��k�A�pr��y��V�zV��HU�m�"�~	q����q�6&3I�fJ3��`�-%���ɤ^�t���3(��rq�JS4���6j*{F�0�p��Ӡ�$��{�#�����s�m�o5Ȅ�����W��k�GB��nѸx����Z��ɝ}��� �9 ��~��;�/~�`�����(:����܅۝qh�u<���tW�Fc�}�M1���Un�;ܠW\���+yC��B����麻b�����H̾	���D������Q��ٳ������t�eI�x��u�)qR��n���?�\���-��ڡCÛsO7����X�D��@ʙ>w�V�>hmU�+-f��\`�s􉳶��F�f"R�����;./��ihd����D�鑰���^���,5@��<t��a��_/ی��Z�R�-2(�A��)\�4;��t��
K���}Ar�&�f����3����2J<��0Ls\B�/q�O��c��^��Ŏ�DO�6�%� (�j
x��V�V> t�<��q�6JH�Z�i��8���E ����Jv����/���b<4��6r̞��}�l�"����t���ʚ�|��?��#;gy���a�V��I���y9_x�]�%�@��t��B���z�W�t%Թ��^'=��� .�?��t��8��NG��#Xq�PXMV�K��>Kf1�H������/A��B��x:]���MM���a>������@\+� K4�f���W'��5e�8��ƃf�\��N�׮��w��
���b>��4�/�?���Y��x�%T!�BE�f�\�U�c�;*ǐ���'���Y��lg�
g�����8�/�@uLuhdw�b�3$u'��az���j�V�J�vj~�D21&�(�l(�+�f�t�(ء�Z����$ �ڻ`]��{�	k-qZ��}:WRD�2�ۡH���Dїʕ�㠘w�WA�G���3���\����8]��{���K�n�f$ƙ���Y���9# ��."�����y0��Z�/���y�Q��=sѲ�)JQ��1�wdVu<�E�t�4K��۠~+�i�~A���8�)�Q���t%ٗ��}	�Ck?�R��ᅙ��F��$�����\.|~)пs��m	���A�DE�r%���~����պ]ŜDl��r?y'��T L�Xh��,~�mo�6k�3&��.m��h���P`8m��E�'���	>	V&T5/����?,�2� ���^�?֍#�f�=h	��o�@Z	���4��H�H]�������Ƙ5���q=9��j�#̕Ow��q*v����b��8�j�d4���')Z6Jc�P)��w��'FJW��9�<Y���H=�4� =�;�{`cH��Pb��'��o���gր*���)�H�`?v�t����Z���tz�4�&�o�.�}�e���^$U�]ۻD��D�:� �u����,6`[f�@U�'h~WQ��o�鼚k�edE�Q*Hf��S��J�=���{l����o,��|@+/��h����-`%9�;ǐ�����QSQ��4�N�'�<�}v��8F�o�e�a�1��?D�ɴ��;.#���/�H�Ӡ����X�f�y��b��8�[��p�M�[>�I��`��T{�#:���'�s��!|�a���Q3uY��h��;��?C����p ��]�;q�)?&�q�}�ɓh��V,��릔�����T't�:Ɛ�38yoa�����Z�P����?u�D����zB4X]��Hn8/��X���ⲃZŤ���C�#��cX����E�R(�/�m�I)A#��׃,����$ݑ��M�g{�6��g4��f����N��ʁ=�������W~��@���0 �	{�%W �\�&eQ�s#OvCQ���3>���F$?&��E���x�_�؎8iJM�٭���n�~��-U>�)H�&{��f��֤�����Y�T��/�̕Oo4�1�>�Ϟ	Ӥ�/(���*HE�LYs̑�����Mf1�$����B��]�Gj�>-g �M��:%�'k�O!�ڌEX�A觌��X<�j�F��m�,f6K�����Y�r���^h.�M�,.Q����Mrؚ�A��G�Ik�Z{-�e|�9�q���1�B21l,m9�R�OctN�a��(��:־@������V��@��T/����؅؂��,?�9s���?�#ءR^���A�ڊΗd���ԖgR'���3#	o+n��'�.߲�g$�҉��m|jP�E��@��v �(�х�P��ߝs�\�i�F��������+g�DL���ʱ�s���.(�
�.+ʎ�$Y��������F�άYd�
�>Z�4��cq-�&6��-?Z	�9mRK ��$m�~���d��	��ua�]��O�}���J�1�Gj��=��{�F��GE���y��j���b1��f��^+����/������ l�F����A'��?�9eɇ�C�݄'�GU���%�e����Tz>����N�=��a�bN�H�'�f���h����WV��VW�]��"0��dËS��Z�k��kGE,c�$�A.��P6\�cJ{P{�7b���r
/�Ң��(��
]%��y.������Z]�0�IM��0P��Ka�}��:
�R�� ���A���g<{��y�~kb<���U�6��2	�h�����IBC.�q��~�JL,c��RY����曑�K����CAI�j�A����Ĵ���R����p�Ģ)�]��(�D������+�fX�3^mzA����?���(G�ky�gR�[iF��Aڧ,3ծG�7��[%6���1��P]Gt�~�=�g b�%�4g ��A���<���Ӹv���a����`I�`��lia&T�
�ᑣ������,���;? Spc
��Z�s��gL�l
)��F��RpR����D
��.�Ly���z�2��>���X/��dA��b^aS� �2�V�>�QG=X�`��PU�W�Ɵ��_f
�OJ�t��=ث�H�ߋKK�~����a!����FtI}�qL!6Y���/�3�5=��2�p���KMz����G��۸��	���"�e��y.]@a\���3��y�.K̮�#O�.��-K�\�;X\�~�I<5� i�q��F�
�1�F�A�I��F��-�R�\��ʙ����u�����R>;���k�};js�Ã���������9��#�1�M,2"��S�=�BͶ��D��s����U�5�R�gt��^��Q�aՇ���lm��N2���`y���o�LA3��p�C�Av��HK.W�Xgv+�oT������<��G;���0�;����{�B=����x	[�F��G�?t� I�)�p[n���ڠ |�ُT�p:����'��>��T&��S��$5�dbnnq��ᠢ�lȫ���
�C�T����oT5*��}�|�*_��z�2x�i��qn�����mq��е��Lc4�zG�dvY��/S}L���"Я��OV���%e٣h�,(��Ip,W�O�
����[����k%I���|����8�����^>��O��U����N��.�T��m ���\�RtWc����A1�c�c0H�K�^c?Y�0��i����Ǌ 2X�u7�qG�quv�9��]���b�{��8�@%50A� u_��G|�ε�7 n)�]Qb%h%I08���!6�d)����4����ygS�g����k�o|	�BW"p�PB�"
�8'M�K`�Cq*��M�b�ٕ���v3���G[/*sS��,�u9*]�W�����AB�b<��E�)����q�`]����4A�2+��9�� �՚R�����~rs���0� p�6�j�����;�R�"���@�in�_=���s�
8�ȄA�W����eY�A����Z�C��)%��R�L2��O��֕�[/�x���}`}IC'�{�侼ԉ\��E��WS���aB�q=��o�N�PM�n؆��l����;x����d|��59d��NS<���+�4���g⛋lXB�1H z�ݠکoނ�����d� ��$v��m��ثD5�Yl�
?�msǵ}w�&�Z�.�~�|s�)!���O�r�A�����wZ=�$�P�M�5I��\xiv4�:�-�M$9�T�,[� �_7����(*`�����z����WJ����ݭ�kv��t��}��cS�M��!�\��y�t�çuB�R�>������/u~��=�>�Ct�8#�Wק��p����E���%���eUKLm��,Ew�
��^�P��.����:i�3���S����m@ �KJ�A���.�����\^���w�=��y�3���I�2�-/N+n��×9�c�C����U��RL�)>{�}d�ѸN�;�R	���V��3$��Zx�NB�ɔ��=f�U��o�y^GU@��� ,�	a�����L�T&��%j�~������,ק&���߈?�v��	Y�S>��GX��1�G)p��+9i�͡��ǰЗ�|����ߓ{�/�	�޴SI��t Sޯ%����&E�p���]�㪇�.䀫��o�ܿ��<�-�2���I=��=Q&,����qaڪ�3]�����,�K������gK��$�{�`MO5<���k��|��Zŗ?���؋|R9�h/�.Ҥu�$��jܩ�֌��Z���f��_�7X^���C��t�Ç7���Zi��c�L���7#i:��;��I.Se/�<�cd���v�:ᮮ%U��u�����{���`hە�l½��3�k����h)˲��]�(K�h.�}��>G��'ap��j]^~kץg�7�����m��?>�GR�t&�ĕq�i����)��E��G�! ƅ|Za�f;�p�c����qХ ]>��+ؿ5����ϻ%����plߘ�|�u�.Z`���%��q�i����e�(�ȅ�������#�<JKC�C��L�L'�4+м��z�
�'�ީ0|N@@ ��^I�61�ۂ�-���㱌�~�ղ{�jZb�_�����z��>���E6x��ܵt�����B���,1�U�L&�#Mzx��%Ut�c H��K�s5_�����=���)�<��`ٍ ��^��8�cA7~$����Ger�*�l[`O��~�� H�K��Q�r:���63��0�I(�Ɂ��v�)S=C��(ݿ5o��g'����%eNZ�Y�Df}���X��ί��~&<ӡV0�+�1W�\���@���A.��+���T���8��фnQ�oa##�s�[q�3��,���*;�Y)�p)��>��&�T��_h�y�gy�bf~L��Ǣ*(��ǎX���~��4�KC!�\ow�-R���u���k�i{��� .�L�"#��@n�dYtq��xr�g��1"��-e�2ԉ������:u�9$���=�jĺ	p���Ov��2�i�������8���=��{�V�C��'5.u���-���o7c�)0K�i0��q6|D�aO�x`��7���]��xD�h%��߆�߿�u�Y_���p��r��T�r ���J��|L��,�8�������o�
\�no��̞A�$��yTTb%��;_���Ƭ ~ �$��P�Y/���b�K0c��9�!	�"y���Y8�Kp^��J�m�����^ۢ���n
���=����z�/}L�Y jX�ְj���t�����!����m>��.þ�߁Z�R@6LR���D>���?)�$_/~�+;��P|��^�#KLj� ��9�qُ��G���6�=5�5�0>�������=��ω �v�-l΂LW }e������0���.���K �%Q��ͨ\��	����ߛ��i��c���`�J<ITcU�����S���Qe��Md�7�e|�̎��-A�J&�xUO��>�˹�9���<ܛd��ג{�0���ߗx�h+��C}'�Ny��,��d��'�3�B=f�u.[�D��o������^
[��;Bc%�&����*ӽc�<?�/���}B�ٷ�P���hu!{�E�5f���oEc���r���*h|�������G;m�5`/�.�����2����汸*�\Ig:�	�"
��*"@��#V�%�vF	ف�H��c=�<{���S�J��P�	"T�T�/|�����6	�CvI��vXDv�*P��#)65~�;�c�1q2��LT~�F�!�@��t:�7m��*I=ˢ��f�}l�����R��WM����	�?82��}'r+~2V�1U�ʑU^����OZ8PCc����_�If��!PE��@5���o�݋�'$G�0%�]X�8���/���U�	c��]���_و�d��?\����&�ҘM��nyK��t����q"Q���J}�h�F�VW�(��C:/q�X���������B�5���0��⏿������
����:�IZ���C�_�[*ˁW%���8�e�����x%�Q�8���� ���D���)�,6U|xR����i�_���a��X��OI#݉���ݫ�4�;����,��/��JbZ'���.�LN�mы�9��4��>�o��7����noR@�b,�2��'���z�VD��' A��"�m�S�}�$զ�*����q�T(�)�g��Y?��,�j�,��tQ��\`I[�2�B�g�m��O'C�:��<} �;1-u���@9v�Z8;�[@�RK�D4���z�H	�
*���?i�ߓn�e�ߦ�2 ͼ��75��u��)��*xEե�:	��[�L�ZۡU|��p�~Q�&"	�8{���dn�)��׼����x�O&d	T=�3dri�TS�Po ��D��)#�ޖ���>���T��:
A�L�/6B��B�9�|��
 v4$��6�+"��6�>�Pa�����~_�$'��Ro^��"�aU�BA�������	�����M�![,Z�J�;�c�:�Ͻƙ3��pa!���;����l"��N�:%��2c/�N:΃�g��n����.:{s���m��{nv��A���t�oK�\���NE���[6{��_?�2l>�XV���q��Ό���YLu�)�1C�	*:�qn7�ĶMzeM�}�KLY!��3���:�v��ŭCYa$L�9���+�(Ք~��b��g&9��2��[m����(i>��-q�,ɫ����G-��(Z�,�i�y��Ӌ�5
�i��r6?��7���WQ��E���n�����69�ǤԚ�j	]9�;p+%� �co�e�q�����<�����g�ߊ�Zң]YX�L�.H>��>�j���g�׃�����:�����UX�[l�{���v��aX�w,��u�hk7�C�J�ՙJ�w3���-�+���B��u���{N�kLgQi�U�J&��g���ku�D쎕i��J��F>���|���4� �Np֘blo⓯#���9$�^ ��{d�.�L��݉Kٶ��,=5����B��
l��(C~�X�[�v�A�$1ll����E����Ƶ����7��(�~�DZ5�����Gy+���G�<��{�>5@o~j��4�wn�{yHQ���y9ቩ�(�'ׂ��@��Iã1&j�gEa�GS�7{�[W���^Oh���O���S�4���eD������"R��x�_I�R*�S!>��(x�u��?�#�����u`��g�;����Vu65�" KwE��4��H��=oǺ.�B!�8|�]@_�Jd�?vk]��tj�d�2�=/8���/��9�
Xů�Q���m����-BQR��Jd���	j�2rh���8��S�t���od��BK>�)��.M��~��VcPȻ^�!����Uכ ����8�~b�$SW�'�i��Xb�B�>�/.l��.G����F�?�~ �g�u\�@�e� �]�cڴ�"󓻯���#!L��B��<�]�L̇-A��-��	%��c/_�Γ�'|���D `�N_��?lnyZ��V�\�G�"��&�����e��*p[EUPc�Y夫��T̅����=���S�>���@%T̊#93Mk�iR'rCO;Ϊ| ��1�����~��c6ƹ�h�"��!@�@�Y�.]I/ɘ�\<�K�/7�J���t܍\�^�^�
��|M����K]�m�n���<
��B�ẏ`D��j�$���*-�M/P���eR����T�JN��oSp�Eh�3u6��E��fբ]��� �ag�v��*I,P��;��T�L/�v�hʖ��v�p�����΃�������1�#6[�a3M���zn�}@-���` �;�}��*���?��y7��oPɨ�M�F�ȸ4�&��fM���ůz��3d�2_�%NJ�Թ�c/#�~��G�����	.^�g�iג�=�TG�l{jzF�/;g�T��6�J.��4�s4?�G��7�������(�� �m�o��z�S��w�%� ��j���@*/k�G}¦��Q�UA�.�#��$�t�E>��Jd�(�ed�r|����k�,�z6�?����ГJ��VF
�n'8��/#��(�&�FfB�W�/2�*����d?(y#I|���d�E�geSkPe�4S�N3�$$`ܝ����k:����,�q�(� :a5������9= &+�����8��b�T�����e��'1k8�5iMB+$b��
�$����f)�!�S�L�4SU��T�߻O�y�V�Z�+ar}��ʸY��c�;����� �ü��Y��1�]�����ȅ�@�vB���\s[���b��lu�����-��`C�M�Yy�e���2Ǭ��JO7\v���+�Ϫ�ܹ0%f���S|�U�w��Yq�>rE�~l�d"�SE�_�0䲻4��џ1�U0�-�w�3��kq5&~ �:9㴔�1�?��������^+��yyD�;����-&֒1ϸ2��hB�lưA��e��I��RE���ҿ��B}��"�f���:$|l4`�%�[h���4���,h/NΚo<e7�x	2�ᙽ�������������Y&JtY.RT�{��*����:��Mr� ����dO���<��``��t`�&a�ƻ+,���3�<x���ԟ�\��o���`0Z�"H/�G�	2��f��{Cpk��Cwz��[�^�c��%Ũ��)�,tTI�m�m!MQ��~���46�ǜd�{y5XX~ȔG<��c���U�֧��ݯ�k|�Uؼ?D�e x^W�D"x-���l�:,N
k��)�0�!�|y�G
	�5O�jK��?�yxT�.�ˑs�O�V���D;���>]4��W� ��F��/��gr�k�n't��y�,���j?T�n:��_������S�m+�ns����K^����,�� r�7�GQ�x�y�I�<6�=��l��x-�p�Ey��y13��7��ݽ�(��L��� ����%q1E�^S��h�w���2,��W������$�硍P0iH(�G���	}9Đ�n݂o�:�<��2�Pm� ���p�KY"��J-l��������g�����Y�Jh����	�w���"�'/&�0.MB���_K$\}�b3��(� 2�O��9��A\�'�m��iC�@���Ly�P����З�1x�i�5�2 ��9�fQ�k4`/Qϐ�l[zH���Zb���a�V:�]<��:tm�����h���!Mu�'�v2��ħ��P놀�*t$!`,��9x��n��"Qtph���߉45�!��G��R?Д�j<ާ_���ɮ�$ �X@ʝت@	�3�_��#x�"���ʎ�� n�x�)~�G��:
�@|׿@�+�cٛ]�\{;��X��1�+h���Ul'H?s��VIfÔ"��L�P]�j���5�������۴6�O�������� ��REy���
i�K+,�OB�$���BwV��g�ǽ�
���?~B�s�@d�i��`��BЎB��Xw?;"5�h,gE�f���:�#ݯ<wX �<�k
��Mn�)��-99=rh��v#�ϫ��,��ZFo��
zMaJc�=lZP���]EĞ,`���h�v��	�������0��2/��R*<ޑ��aD%:�u�E �ZK+�;l%Qqe�y��K��Ze���Ʉv��%_w�Q��C��a5�4 �ǐ��į���k�e�b��S�9����Y.��Q��t�^ V贕[*ĔW~TJ���ۍ�9�����Ͷ��`K8�I#z���󭈐)( �ӽ�}O�=���'����Z���`�%�^g����R��L�`��KHpd9-"���A=�ݹ=�x���3���?#�������C����htb��x�꽂����^B�S�ˣ�U���q���t>�־��WwX��qv�hy�9��pc��j,�΢�[����&��g&e��]2�jÔ����t/���䈻�u���Ȭ��no�v
�^x1����*O�:$w|�W�]�l4�h�p���_8[�$�2��:�o$��1�i��,�t�f'�o �`����p��g�������-����{�ĥ��p�j	^ʬ�~ �0�L���c�\jo�3�#�aM����O���:�q�J�{<��.'q�$XQ��Ľ���XHY=��抂(N�n|��xմ���Ҁ4���mj�>Y6aɹ���> ��j�'8m��|�G�PD��
��r���FU��Ȓ3ۥ 3�����l��q�4���@���L�� T�k���ϵv�"�s�Q��6`�_��Myn�����;�1���%��@��vI�H���V��y���!�.�6���;n7���q���>�2Z��Dw��x�Y���#Eہt�#X�(���{*��;~���<�����Uq����8�ӻ����� Gd,���$h j��F�yl2VK�>�7�t
㷇��\�gW�M*�t�}��r*ClէC�{�S��\�Tc@b�=x��t�jc>V3���/�b �1�v�x��;(�e�d0(n0���d�C�u��z��GD\�J)���X2�-y^�A��?i��y�5K��X'v�=2��Qb'��_ˁ!o=�v�$������*�l�z��ŉ��V�Pm徤�����y�u�O<K���P�|�o��拁�m����ի���yyc	�2����q�Nz]v��A�J�'�d�뛮��QJBp--���*(ָJ��O�P��|;ri�����{.�u�C�����Y]�t	���cW�o9X���P�}�_���,���~/ % ���t[
3*ԋ	�Y�/��7XQ(�T]O%���A3.7���!�iBy~CG�<j�bH���͞��v-�,z�l�&cJ��S� ���)&��z��
}���c^{�Xc�Ɠ�z��W�5U�;�m���{nKW�,:��b�>P �s��J�&�7����XOB-(�`)�:��Vn�\O�9�){zU�n�j΁l&>v�:?>^���9d}�=��B^�Lvl�7��\�.�6" �=�C� ���ڡ�pC0�rg��@~�v��]�q����Mn��Da)yO���K��%ls�(��V6A-�0y���rH���[@�>q�;VM��<��
�)������5�Q�IqؗS�S1�b/�/�m�����]z���|��ϧ&��اsG=E���T�5�x�	.�lp蝵�0���Caؘ�o�P�z��e�M�ke�u����/�&s@��di̍Jg3YCܠ)__���̻L4��RQ?Ɇ���$M�e��v�91u�/
GG��J{7�	9sQ��?!�2�RZ)�tň�����|��oy&?�g������?��,�cn�^��d��:���Rj�ڎX��D�p���~�x2�%�T�ѿ�3������er]�S�z�~;�hE#����I̡0;l"|"�H��£kQ�_�e�������w�#p�?A����XN��w�G+圫���ͅ���H�R�q�*&|�5��`\�*�k��Y]�/��gܵ�	B��S�l���� ����&�(��i��9�Q��tp7`9l�"2TC-B�C�#����I�o}P���eD*�t�"P�R�.5�m�h9�u�g�V���E?�p-U�����^�h� �t�ʬ�=�"������ ne[sP�{��l�?U������o�OT+�1�NHE@�* �����j���ϸx�77b�	G\��Ve���|�gf��
�N�P��^j}ZAu6�T��#�W?�c�O����&@?�!�M��[��¾/3�w~%&�jEVamƜ	u�o��;��� ��q��v��,���Ӱ�v\'X��]�-�J�
'n4e8���y�^yG�q�Ɲ���'ı�A���zǑ�_�6Q�W�9d1��d�)m���q���j���� ã/��ڮ��}�.�J�׿�(-:`���BR�y�h�P�E!��6����Q����-WC!���2��|�b��$~�(�y�xz��|���\����1���e,�݄Y%�5�}���yQ!����C�������㜇�Lq}�0��_Ta�Ot���xg8ߨ ���O?��҈�`��-�}��"�C�.x^�(�9�-��rm<Bh�W���zАjCJPd��U*)Sʥ��8��4k_w�$IA�Gh?U������|�:�P�.�p��[u�����GJ L�?�x.��&�շpFG>&8�M���G�ar�������s����R�N�Ub�M��'�myB�v�6��]E۳�G�s��  2Q�4^�����X+k�������c���V��+���7wO�+@�ݵE0��%��y˹��̰'��7��c5��j���n��}�L~�ꕐJ�n59W<h�gD���M����}Ô��:��O���jq*�aa���C�E�c���2�*��QD�Es��nw=�R��,�6�h���r��f�ż'wW<p���`��X7 t�ڗѼ����v��j4�.k���s�;�|��F�"�krg�+a�B�U��9��}�	��� q1�;����*�r1x@s:��$<�C�	{Q�}O���m������uS"J���B6�����7��R�H��Z1���	M��5��F�} j��J�I�*2���xSb{��|�	�#۫��Y����օ�T`C�ܝ�1�s��z����cx�R�g�6,��~sagqJ����0k5��r�zj����(]D���^���D�@�"�B�Z�n��� �;�?��Pʯ��c�^��Z��[�/Dd�e�i�{QƂ�<F�Y  �|Xg���t�#�z�bF����K�N��L�t��c�o�<�y��{�ϙׄ��������̍`�a+�c��D�`]ҁ[ɿ����	q�p9Ӆ@���v>��*���v��F'/���bW~��Zmy�F�F�)�Z���1��R�Ek��E�3� �
7��[��Pj.�\��E4T�%>��a�c��o�6x�zA���%��2��D�:��d�@��zp;��c����	^�j�f�;$�ـ�N�2�e;��?���
H=�|q��׶�����{�~�lpz�}?��s��d��HpA���a/�]8��H��`�
�z�s0<��*����O.ňX>R�@�K!�D�n�ǎ�
ݭ{>`�5��}����gl��oAu�q^\?��p�w0G��n��YP��_��:��2ǨBu6xe?��]u�ͽ~�7��� UeL��R���g�};Pܮ�V7���֭�i%��&���T���4)a�N*>\nʗ9`��S(\�)lV&�Ə@������� ��9������抁,Y����i��ߑ�X�H��x8&���Խ�	�$g)�k��|����Y)�1mr>��W���z��Gp9>���Jk�*L<^�U�m �3d ae<I�#ٹb�$߄��A���En�l�ցi2�⢬�,}$�DĞRw�m�y�1�W��D�A�y�">�	�����×��V�b�rP���ɏ~'˟�;���TPx�7��	pڪ�>Wϖ�H�v�!����A�cq[���ig��'}��'����{�>�S~ЏҌ�`�:;��PC�uyݫ�Y6�a�O��R��L"2#��!4���~#A��T���ݝܹ��)O��) A\1���#��O"��u��XF��j��ܠ�j�Ѩ�&��op^���C���UM�mT�i���G��{z��T�cm����YoxBA��9u�W_Ҩ�����A؂$�����n
7���D��9�6QG8x���!l7�t�����t!�@�=���f�:�Q��g$��9�
 �pK A4�$7�H��F��4��FsV*
k�T���Cu�̐��w|)�6�����rAo�����s���;{�9_�1���y\P)Z��R��Y,'&W.���JW8ϟ�ק�)�V8\�'��F�̺�
��g5�O��\��,ӥ[�Q�q>eQr#_)g1k�|	�� ����>{,]3,@v��Do�%�����%���k�!�%Y!tI��1��R6�x�놪�y �,mӉkwj���7E�-���L�shK��]�X��� H�Z&�ӄ��_h��
��<�h��p�.TL@�.�'�ߎr�f�o�}��15<�zDs��?+�8�҂0����]-���TƸK�ٕA��0�gIq�?�G�9)|�u�]Lm\W/[=�3aky��fm�rs^W���-=XM�ӄ�Gf�':����L	ɀ��"s��l�r�p����"[A���D���U�@GO���u�]֔�`��->~�2�W��X����n�Ȁ`�F8\k���Ķ<�<�%���7r�p<�eSH'KL�5�b�TN:��e�ӑ� �9�G���[����tJ+��"�T��9Rc�C��,uD���Y`�"��&�ڏ�x]S RuG��P����	jY��6�F�-L&�.p�&�ь:�hd_����:5���*�͝$;຺8䙩��ƎeE��R۳&y'�a�{8������k)��o,�;`� ���Q��V)�Z��"�$�hd�U:@t�)�O]@�U'5��\����A����_W79m���<�P|��W7�I���,b�uE�R���<��K,�ꕶ��>�V3gcW��)[F�1~�&Q<a.Ne8M����4�B��ڪ=���~��z�]�`S�?�3�� �H8�E�-��2EĦ�O�.Ȉ	zS`��3����3��N��]�of���;F9m0b@CF�T]]�b����Q�'���;9Ye┸+@�;ܾ#�/6C�L����+����G1�jS
�KIP���	���Z�"w�9�{t]'�����>0
�$���,;��'u��E��#­�<�H���R�����z�i���,��pũj�10ĵ�X�����fp%�ڇ���`UG��_��Jv$�
L�ý��s{[�^����cB�Y�c��{.�c�I;,�Nc���*�A��D9�E8�S���ǒ �W����D��uqs5m��[�Eg�GI��n��
?�Ǧ�|��L�y��K�2.]��ӎ��<�3<��$U��lu�K)z"O24?.`c�����^����W	��bm���mG��҈�꾹o��;�7��R���R?�����S*>���Ì��D��j�qK��M�_')uF��*:���8��6T�#�5!y��&�*��]�>PM?�!����S���	��;��y��i�x��	��k�؉�v��ن�6���hF�<l���P�����W��#�[�V�3%o����>Z5��&����j� ���N�}2�C����1ƭ[�1#���N�K/���������,�s�c������N���HѰ�Wv$A]��7M§���\�}�G�s���Ƭ��!;���W�Ku~�Kj� %��i�1�BT{e��$'i���L�NH=l(J��S@�,PY�!�����o����S�۳J>v[�<��=:W�%Ly*J�/%^JK_j�!
�[n͍���v�)R.nh��?�z]�2�o?h+h����d�;�P?f�����
Q]M�H�3s�c�vXlSΣ�f�xچe3��9�jz�0��7���������d��Q��y��@�c���OI/�Y<pu���2= Y*�R��5m��ޟ7�� ̾�I|��Dv�����AՃɼ�D~ՙ���	ꄽ������@��F��!.n��o��nf9�	�j��Ѩdn����q������C(Z1���~B@�c�����h�h}ν�q��m��Ǿ���DB�6��gv�/�5E?Ύ,1ٸ���n~Xq,Qoaw�M/P���*9�a���DI/�Џna����Uc�,��% �CN##���T�Rn��0��ͦ�sA�R�H�cg����.(��]+��#�l[%J<u�:_A�c��%�4q��O;+e�����PQXh�*uG�����#ZGw�dj��Y'n�A�_�������.����W:|N�?��fI��� 0]��R�#)( ��	�k��~�A�� (�S������v�!����G�%*,�ܾ��L�4_�i+��d6�Oda5���Ab�!�J{�g~{PۘՆ����$â�a��M�$=|i�v�b�-QG����Ղ��b����Hړ�߳���f��2$!�p�󓸸��rZ�P��3�k(M=��K&�-�<G��kk�ӫ�m��y����!����� ��X�z���xu���<�j]n�TO��	@Pa���(6��p$�H�Fs6Wjԙ���z���͋�o���n��:��>�WI��F5ܮM=,��kZ��]��kŞ�h�T.�[���>S)6�d�D��ET�%��#4�y#��Bx��$�H�m_L���zw/	9�ҷ4|���k�>�NN��q)C��=c�wl�����|9�.���נ䘌�kj�d��j�ԕՄ�^��q%��f^���M(����eőDGn�<����_�?���-�o���a�)v{�>7yi���QtO�G�.&D��
�d0|2�l� �b�G����6RM_P:�T3^�XW
�Մ�<9�~��(�%�a�M�y�$�rAFs+����n� �8	j�g&���#�Nb@�B�.�\�J��_���;�U$�����3��}�S�iЪ�Lڞ�-�����j��
�5�f҃`�n��ݥ�iN�����F��<����"����v.ߟ�T��\
GX���{2�w�1]�Խ�u �LO��"ō�'_@����M|�";3U<��r�/CB	�)��<><!��Ү�M&��n���L��f��kQ��q�4H&!��Wh�HY&��uj�e|�#�ROb�  n�<qc%�9��'\�xJ���i��c����I����=���P՗l��C��� ��hb�AtR^����B�V]�X/Z�6a�o�,���V*����1}³l�#d�+��0k�ɞX$�*����G��z�|h�u��Z����B�����LӪU+�9 a�mu��C��.y���I�%-5<t+3K�INFZ�9�G�(r;���ݒ,����I�����BA#�k���y�RF}A	d��r���IK�,���Q�26�����޳PH+��� �$j��Kc~�`�;m�A����tn���,�:��+;*̌ ��fL�C���[P�M�`�?�AO�֖3Rq"`5b.u=x���^=������=��*eyy}��*��Y]C�Ŵ_��6�8"�����@�W�a��n�z�$h��V&Z��j@!��	�M�X~0��~�P�5r�$j��z-ӫ�ɺ���*�b���`��0���x��Όs��뼕s�cf.?�ÁH�;�S�%;�|"^p�������@z��4!cnӞk�����ͫ�v��#K�'\��A�A.��ԤbvL�-�I ��?�>�As/���쬃8��pQ����% J�aU��H�טc١><p$��y�Uor��>�9�l��mv�W��(�s�v� ��F��r����b*P�_K~tq�@{pޗ�D���c�~�f�}��Z�=�C»x���^~�k |����x��/����Kc�]�F��oX~1GM�Y���-'~y,��\i��GXj�z`d�'޿D�	��2,��N>l�.&���3�'� �di�R3_2�%q �t(J�$���=��]޵:p��#��{=2�|�/S����ٹ��O�f=wm�LV�s�&��[�D0QO��Ta%�@�.T�4�w]�������ƔuI��^��`	duў��w���a���?�-Q��r����n4�):h�6���J�{��L�v��]��mM'���e(`��!�c�PYs��I-��� ��g�4�o�U�O�53`�,�G���4�j��:����ym4��q��V��+E�d�?�� �C��B���a!��$��ӻ^T��M�/��=�p'�H^��K�R��g�yz��ʦ"<�����c�!9<��\��C���՚<����Y��нt���%9��FG\C6>���7`(N�j���-o~`�$�Ge�j����F���~_�ь�d(���k�_���%]\e�k�\R��#h�K����ۡo$��ͮ�@Z�����e�]���6�ԏ�2��āر�V���/�k5�?t �K�z�F��L&G��>�a�[:��O�m���M��OZJonDK=��k�*��\P��F��8�f <9B�m �if��h,8R��I��ߔ��4�W5GIjV�۲B��=ų�>`�5���嵓UhE���1.t�DOjd�􋐷{!>I����fl��5ӑ��'�WC�Vuh���;*.m�7��W�:��� u�U8?������WN��3EHS�*�;K��q�1GWD;}��3�r?�����)��a������6.~�����J����̉s�Ȍ�u�t����L���Si ml�?�������*Q+�q��WY���<�0��r~�5��z�럈6�z�@k�v��cXwn+��:��?��ލ����l��,��.��y��9*yP�3wi�~�L�'���`��[��6�T�9�VJ�K�h3��O�)W�<�x$�9�Y�$�(-GM#H�J�Ńwm#��4��jqe�'哷H|��� �)f��i��*���d�*�*(�6�U�*_Gí�_]���C7�Xr������C�X�ք���p��+�H�W~i���O��c.����!h�{�aj�� ��!��0�I���S�}qE8�F{��L��[B��9%�����2�k���l�v���>������Bb����3��+���t�� �D)|Q�nxR�,����c��U�(i#��n-\3n��XFlɀy�ރup���a?�Uc�ٻ)�]��^����Km����m��0n(1�
�6���7�\#�Z�4;r���NK����NM�SҼ?���9���ȱ|�(�K�2�^�(�'�E!H�*��Ҙ�:&�����M�tD����W�ڊQL]��zZwM�|؜H䫥s��E�����a��Ҫ��[����6��\iO�^�I�Vl�T�?��;�U�+��4>����F܋a��ڍtU;p6�'n��F���)<0,x���{)k�Π{t��B0,�[��-x\(w��e1�+T�f�AK%��$���5��qk���s--dV��&y����M\|b�����!%�z�J�؇�L��?�_�@��U�G�sNU�\�JE+��Pü�(�����/os��F�͛r���_n�0=٢%� �e���eM��2fj�hn����V�"����hwg�ʴ5��tcp�绠幼z���@ؒ���G�מͷ~�V��u`=�:TM��)Ez�l�D�qr�(��I�m�ee�;)erpb�����V�%�����Z�=;6�]��Ƭ*|�o5��o��h��Uw��f2�/��W�Xޒ-����DW��0����tg*�_b3�T��AС�$���&
��1�v�c�H��9���4���Dvm�Z����!��>_�k�H�0u�B��VR��@�L/���F	y�p�*
u{�,	3��ˣq�<��^��B���Lx�_��EIo��&���r� $:nfVXrͽ���iU���D�8;=���g�^_���1�2-)2M0�Ӵ;�T���~����G=#�����0!GSM��Ld~����K{3��5	�.[�N5����tW�a���ߥ�&H*tñ]%�F%5$	CDu�c揪Z�=�g�HЛ��WX7���R����y�6�BX����H�қ_13'�m�~P���z������H�ݎ��uSz���7�S���`��Po���>��l�5����V+8d�^�A֦�N0Ik�s�t?e�}�D�� ���q����kU�Q�E<�0 �n3�S��� 0��[�ix	��⬫�����n���2�U �ʜ�t� ^.wz�yx�x� ���bZ��Aǉ������j�i�U<jNk"cD�Eo����˓K�~����r��O�5=�4U�r`<��m2�Y�h���C�`��G��nӚ�E�5v��)o�F�;��p�UYb�E��u}{�p�U�����	8����u�
wS\" �e6����Za�P\��rs6'i���J6ɶ�_-�^iwk����m7FܼYK��QWѨ��^�g�F��)ɸ�C�� 3�#���v}���[�8;���k*6��}��K��5[�����ބ	��u$�>C��������cr0yFڈX��ƽ\�G�lb��;�8�w#$v�­m�s�&壟�R��rw�Xt��`��%xf��pEI����-�����Q&�t(1�����gq�ފ�I��\Q��`�!�hB/�J�Z%~�$���26��g��,H���IuH�,�&p�b_�[']%Qa����/C�<�'�d	�Dܖ��K(3�>�f%�Y�ι%����s3�9��pQ�-6�D�@���
�"�9�b��nۡd%���;��E��Ǯ�am��˚d�S�Ȩ�X��ڟ�*f�T��AC�M˖����}-�"U6�����C��Tf=ZqrΎJ��o?^�Z��' �_��6�PO'{��D��Ww�4����h��/!Gˋ��n��j�q������\���,FUvs�m�1-~�.�A��8-���������Og�'�H&/\󧚳��AN���7�4���3�o��a�I2�7Z���޿V�tC��ۼ6C�
��#����$��(�:9�fb��P�uB꺭؀�9f����	���ra^�,q0�|�I���n�whU7[���7R]�b��a���/�֜,����W
��e�E��M�Ѿ	"r������/�-�D���������"�8k��-�[���˵�Pv��#��}F0Uj��O�q� nY'�v"�J���T��s����,u,Y�r5���;`D�i+�㣘.;>ȶ��| B�{C�FM��ݜ��b_��s`�- �_��v�k����.oU
�-_'��C�4��#��"`uVv�]�1��_�M��d�)438��
ʓz��?a��DU��
PJ5湯��xy��l46<j�kU%2q6��Ъ����[p���w�k�����m@r?���yk���JF8��Ӊ����9L�Ph��D~A��ݤD��^�Eo��+�0֗�L���MC��_~NB/�愈h��?��+�$b\`��*�_`Z%_p���Vg��� �;�m�"���E̫җ_,���Y��,��ɻ�]��%�#��?��9C1��>�����a?�W��{��9Њ�u�W��)�]����s���/pj��\z����"�V�
�m��\�
3i�	�o���D�jG7�2򤿧-Xf+��j�$h���	��Q�p2�~�¥(�<uq����n�"�C�rʟh�=⑩}?�L��s0�
�o�m9m��$�_���&�Vi92�J<���Z�O_�C� ���ߘ-�(�%�2�d�Vd����m�!�
�����}@�k6�*�uM��9�H��/�}�[��ץ�B$$��@��e����3���d&�j��/ l�/L��b�D{k��^;8t#��F���]��U�^��&V�����l�{��_����5���X�c�,�V��:�t�kҒG$Y��I3 ��"�%~�@�ב"9��מ�Z�1GW�{X�W��`O��_8$,��c���}�x*�Y� �A{>`=�3�<L�q�2�&��[;���6Ñ��l/��`Ifs�[��D����6�o)=�����aGN�^q���d�F�r��$"(�y��/9��柄 �#]�+�[�;�vqll�)F4$Si����&E�C��:x'O�^���.���*�nk�i�꒰K8��.�a4���M�22�<d��$m�^-�&�u9D�si�,�Ƈ���<B>��r�E��"#��E�˳ۦ�����X��ﯪ8 JZ�XKVAr9 S��-�O$)�/mi3K��`�wc&��Q�
B�\y�i��P>%q
뙄ͣ���9!��2�
�
5C"����j��D��N"+]��EWhr�02SbY���5�.u@��éE0}y�a:��]���v�]]�z+��}9��^���X��"Uo̊�}��m�+~�_Pۆ����g�����d�|,
�Nc� ��{�G{�j�#(_�+�+�m�����r����-��!�#$��˿|6��,=�JH
�z�#�1[�9��v�������[9/��_x9�����p���qIA���>�m�tM>5-yxE�<7n��2��CŊƋ�s[bs�QG��혝�D���t��<��B� q7�������:��K��Oc���5n%�w2z���61�}2�?۱��.��3����κJ�BU���NYn�5��;�D���j2X��E�oK�tE0m߈k`m,��Vk�5�ؗ0��:з�4��Duz��1�-��AM^�$��`�w ��"Yf��D��:���Ę�zhS��y�,���7Y��?�h).�ڛȱC1�xF�O���,f��#D}
2���_��Xa�������sQ���c���?'��>��M��������L�yi��a?�I�T7�	`���Sg>�Y����!o��wQ�M/K><�8 ��*Io0]��(y�,k��+b�\op:��s�]8�k&��W)(��h/��u�����
���D��<���G��m槨�O���g-ۖ�͉�%s���i�?�B�`�Af�R�)��n-7Y���r�S���A
;nYۗ�j�Z���Y+�d�@'#����h�3��KT~r�����h/�d吳������2�	��+wB/lql�(d׎���Xh!����Ο6(�d�m%��!�Y���?�	i�$�g6����d�K/�4誓�[��T�ݚ�. <l��y�<��*�"��bO���J�����E;�ud��["��PcU���[�'T/\C�S�1���*%�I���l���|�O HU���}��m1����T%�2��
<�bb�M��V~yp��i;�����1[@����,Y4�����s���Q�˾��7$��S���N���i���U�sC����8��-��=zo��맵���YF��m�š��L���F�~�yA��Qo�����J���g�Ae��� Ȓq��|&r�6������Ly��:x�rv�'��M�%I2eA)^��'���t��m��]|Cjh�EZ�S�Q86a�Oy1�De�D�A���kߞɰ��hĴ!�N�]��r�0[�zG	׺N�`� ��@���{;m),ERnЭ[���h�׶1r~{}Z��]ڲ����U�ґ�p	�n$졑}`����	��%G��w^�B��5򝺻��t��BJ���\HgF	"�;����.��<!TCl�P���Vj���/����x����i�P��ƷƩ6^����)|J\�/au�;��<&i�س��6:f>i���+)��I$l��k�&�&g�N5�m�����ց����t����ot���&���+�KN�"\�=h}���$��
9�C�kI	Ԥ�䐴3�� ���7K%/x�DM�djƞ�Z!�5w�22���"�wR	3��_�,�u�?��ϔ��%���-*� �W��0h���򴚌u?�����*�%����1��8� ��י�TH���M&Z@w�B,�?O���9��y��ֺ���K�I�V6>M�����w0�?)���<z�k�_ɹz���k��q������`�R<�@%�b8j���(%��[*0�wp�R�|ڙ��ܬH�O�+D�uW�\�OJ|MgJ�txd+a.��9+�&�\�X�W���;.G6Yw��/���;������4]��,=����c�Q����<�QP�=�Kc+��"��1�� �k�ִ��HB�w���F�c4a�����}�:v�t��,&5utc�+XR�!�Z�.*o�p�����N�s5B[�OoLM"�"�b	���*l^i�5eǁ��������o�[�vV�V�)�1�	 "��uW�}�p�J��O] �N)-����B��XBlG[H	�����G���u����r���	%��,�yN��e0��8��������BC���a����Hޣ�ba���{��]���re��?iS>��e�El����)������B>Ud�}�:�37�-��?��W4��=-ͪ��\KC�vy�}�������Ǌ6_�U����	J�eW���\6=�b�z��>�"ad?K�����J�o3�Y��'b��Sm���@�r�$���jl���~>|���n�ܬ�-�{1c�V���N7v�KDRD� 6�D��^��e�V6�X����x���6����aٷ�,�����(��6�����v�� ,&οY�%�*;$,5�6����y��F-�[�7�$5A���kV�̡)@΄��r8����a��~���H���K���*${�Z7�čp(>�˧��4ܚmC2�9P������2���K�q���Q\��E<��I�����bc��k1� �iy��kyh��.�ujB)0�|�|L5�e^���c�\S�ު�{J�� ��	�|&5�z1'Q�"����z�<C���T�-T\�!s(8/���9��LjBd�oM������~��*5�bB¢i�G�v.o�'s�ri���oS��d���EC�KId@.���。f�����M�J&�Z?=P�+B�\�S�}�:x-��
V#��\w�&�����|&��fl9�V�����
A�W�F�'��hW�+��e��N���m?���A�t�NnP5FR��ȤQ��2$T�R�-��,�j0��茊��vu��6q��7m��j�c��^&\��,7P��6j[ZuB��������V��]��G��u���mp!̹&���Maڟ
�"Y�����&�=�ꎙt�]�W��v��4q7��A�惟���Y���)j ۻ��h硲|�R�RMm�RTWܠ$�0j2G��d@�Q�(h-��C@���Wbatb�]���S��XU/��Z=�b���/�4���,gi�Q�*�E%����	\[��u�/
�{ftݳ^�^�a9��\;#�����h��!L�H���޸�Z]�i����Aӄ��s���I:��Oo;GE*��1gV�X��J��3��c,`�I*r�.i����}�HE�|Ώ�Y։s��`u�d0B��6�b'ޏcsq��Vԍ���$���)���%���!s��C��"��@V0����V���4�<��Ɗ!M��֪�j.�'�T�d��������1���A��z�/� j� qu��6������$�ۖ�
��2P��)0# K��8���V!�{�!�D�1��EWe���#3�����AM����oD��//����hѐ���=������/��{W�q���v���m��+�jH���3;F��H���'.�U3��UD��k4��.�J���G4{[1����Ui�V�/v�RG3��u�^Z���1M�N�2�kx0�Ѷ��G�17��pb��Y�n����� ��/��F�S���Տ�����ؗ�KŃ�t@L������I�bG�#����~ZC��\ef��;�O:RF����,�9ݝ�ֲ"�1���:xMF48o���:�b�?����ᝣI��m���"�
�(��B���}UoO�6��T���e9|��υ��&�<9�`1���J��?�?J��T�3�냴�*���7�������˴̢��V��8b�?,_ea�� g�(��C�P�3����RyV�*��
L7否[�E�K[�mR�����w;)<����F�Ry�1�膉�?� KA/qmn&d�������ᡫ��K�r�t0{���>� ��ef�T���ҕ;�-�ȑ�������V�l1Bz���F�]����Vv5ϦI����7���j�ToOg�B���E~��M��9�绩��I�����p�~9�w�����e.,䏖�O�m������.>?���[�y�SF��\$b�xGS���@O<G��i}w�K����é����I{-�<�'�^r��V�fm��'���٪d2p�L���yx�ɗ&'&(�0������`Tz��&���Iе�:�^m�{�j+�}��ӆHX��{��Жc���l����jB��N$��d8)y&�1�%�B�+](6��%Ka#�Ɋ-)�/����>[���O����Z��`D_ݾ��j.;��4��R����5��NW��TpR�cb\ s̆_�2*�Y��}l��eR��F�����L>ھ�p��>����r�:�Tt��a�$�\�zWPF&瀤Rs��[��oc��+�ߘ��Mڸ�~|'�h�&��9���y���-��9��4�����J�,l|���ۓt��:���l��ޤ{f_���%*�f| uW(T����\G��鷢�vt�����%O
|E-�E�C}��ә��Ӫ�ey�<T��t�X�H�0o�nf'1������u�$[��#��kY�©�Ն	��%��ڝ��ҟ	�)B�	0Z��F�'낸�v��k0�¤n� �S�1
�"�nf�%� מ�]������F_3@|Mj:�x�5����)ʡ49]�R�ڞ��+��rge�k���-BK�l��G��Y�ĕ ��z�����5���s�Ea���_�-t�gD�`�<�e�`�p��mD�LNŴ�N�'l�
�&�変�����Y��lro�a����b���>_�X�'�}z$5�m��\B��~�A���Fz���c�i��%A	�w�}�����u���"0+\
��!�,?o��P�C�]f�X��e��<+)Bo0�<j�F��j�+!�u�>I*�ӝ|�Ie�+�����hF�ʶ�4R�@���r2�gw�Kx>h��~��'ޣM��Ȭ����xK�n��L�[�t��ˁeDYh<�P�f�^�z�#�{]�V &�&���ð��%'��aEW0@Y����^�� F|4Z�֥���"Pz�ߛ$�Զ�C �7M�ɫ[y�a�
o�-I��1Nخk� �X���[�;a��n��F�N����62�R��l�(��h�}�L�T�腕�+��K�`�uDp^5�)J���ѱ�<�ÒG���Q5�g�^�7[��n�?LWATw�f]S��;���L.���c/`F�y�~�\�E�=r�
���{A������#7�Q&��x�!"n,%�?���'�Nq���5 �۸�Ǆ@�Xgq�c���p�̡X�)Z�6'Zg�Ɋ�_x���<,���v�N�d8i�(�&�J�ҖM�J�B�a�d.�i��<[V�5;ՋD�pf��z4A¹[�B��� ��&��bC9G�3J껁�k�
�߅l���ԟ�w�M�ʳ�[ƣs��=�=��b�U,'sC{��n���I�G�i�� f{�m�H�r�;�sLCz�2>
:��P �e����ԙ��ƻ�p�E�8�2�BbY=Ł^ůb	�U4�M_��N�(e%	�\�D-��v�ɫ+��syj;y�#cZ�ƭ��V�ښ(�-@t�pS�V�2��Ak]��H�zN��ȣ�P���UQ���\Wx��" ���������R�Q�7��s���Ip��'��&8�����p�}�.��h�zX��c-�d
���s��Z���`�-.I*�\�Dt!���P�gi���3~�"�z�����U�1�M��4�s��w���'!M5!�\���^gU	�z��'�bPрN���r�Z�q�������&��bP�/Xff�y���]��Klc{)^�*��rv�T�~�Rd� �'�����{'�Ơ��d�I51�e#��>�CE�,�À5:i(�Xf�>(^_F�tj���aqL���={H�~�}'[U^�G5t�H�/�hd��;��G��)1B�(�z31U����bI��+�{\��ԯ�(c��՘���,���E�����$�,F__}�(��eM���7d��Q���d��삑
g;�>iR�tޔ�G��=�e�UM���t�ʆ�Y������b:�����]��I������$���̹/�Fne��gT�:(���\,��8gy�%XH��54}�4�3�;c�N�YQٽ��3��%O���o3EK�!今� L�rz�_���9��@cx��l�7�9�+W��[0QyS/����M<����|q���|��!p�HL���n"S�B_L0���w�q��k{��;�t�5"��@`�B������Gq����?�P��X$��۳5��P.-�������N��0�_M�U�d�c G�I��7]���?�I���0��ѭ�sb.xa��C�
43<�+^|��o�usj�NC�E���)���Z��m*>z�?R�Jt
2�0����y������AKE�'ϋ�������H�Ȥ?��<4kH_'�""�?��%ʞ��rpI��#�qKZs|�`6�}�Ͷ��JD�)�c/i
��'^5�*�a��8��N�^/Q[r�g3]j����-���m����֡S9�+�rE��@�RƤv?�	�jw��vWJ��g0����ׇ��R)hTr����n"Sj?�5��7�/�ޒ��(r��\�T�����W�cR�����8�9���dv�p���;���HYŢ"��}Fê�+`�J>[�hǷ�T�!���������x� b���-/��;����}O���V��sZ`�`P�E{�[���:h\)i6���`~�ղ��u��#[�R�}y���jܚ�gG�T�[O����s��D��*w�L2��vr��J�#$<��f��:�^�p���bJ�S��Y�B�˨��Yk@(ỳ%�8������1����(�/U���ϺfԊ�;I�ҽ�T'?�o���v��k��mBC7�����I�f��U�zT�̝]��p�R�����R,��" >�×���oڥ�ǒ���q�E@���L%�P]��Y�&�9&	�p"!�B�o���cGг�;#�u� �N�Dŀ�� �o2�'�&��`��G>jˍ��"��ml�f4�5}t�\c����_�Q�H""Ŏ� 1Dk����"�7��y�)���5����ޮ��5���Kӂ�&��.9[�x����b����-;�Aqq�K�Thj�nQPf�G��l
	����8$����o�o�$,yY1�_]6\�[C��iL�詍��������6P��&�Qj�i_>P:�X{�Z0H4�� �
W�[-8�iގ�&�p�'P������9zu�h�
37����:�,���-tT�V�ԧ�m����Ѕ�]�pqx_�|(��4PV����Z�z�ۭ��}����P`��҃~O�h���4��@�yR�l�^�nǔ�޼)�|��J� �<�֘��aqOr����}&I�
�+����w�j;�5���ȡ�W��Xxe��B8��U�u����ߣ�&�/?)g�Qe�����uc�x�� ��$�f?�m�#m3�E�����锗	�<���G�~��LC_Ǽ�$�?֘��M�y��nR�;���@(2���� F�J?������r����J�I�@j�.�	�&����@�����Ǿ�1�J.g�~�Y�Ϳ�c��\ꦹF4�Z������\j+$�%�P�9��x�sp��!(Z�@�<�{����[O0���T)�zT>c��Z"�;Oe���E4�(r�ux�_eJ�д�����6ߥB���'c}̚�:�;�1���8�<�J`�mư��\~M4��#EE���[?��2�p�O�H�`�x�����ƽ��YΟd��D�%�vl�*,{$,�]�3p�]J�n
���B4l��}ҏ�^�j��Z������C�9�,�XQ�Az��PU��͖�D7�����w\\������&�.[Û��+F���(�z}�ŭ6����������	�*�CiP'WH�@8#��t݀vˑٌ�(�%Z��.+��@�=�������lK�&���vr/k�,l�5
:~{�"�b*й��b�#�xaԘ�ɕ�U���V���L��,�p�_T}������k;�1�BE`�Js{�F�#5�UKw[��,�à!�� ��ׁ�ƀ�+OT͘i���X�L_��I:.4�0����Y�nU��U�WEl(���dŵo��a�� ��x��f�`\�ڼܟ�?�hq]ڞ�"�H��ɕ�m��H5��"|?_(�9�,��qE�9��x��};�d��8S[[4(�[��n!�1�9�<��\vl�U1���k���\.* xC{��흟=��bW^�
��Mp����w=n,U��9�� {���h-�F�^ִ�W��z4�^A�B�d{���p:j
��r�O�k�� d�H�0�2���	bs�_""�(U����l�W�D�G�Ie=/6�N�����ɼ�ٰƧ2���l��}�6�5`���c)ەlK�c�:�	�:ie���W��`�^ˣj ���y�7�09�1朹�V��X�0���b�~�f�y�RAG�*�i�}�\mJG]��}$i��J���[���>O�&�4ܹ>�x���9���V�<!�\�(/,|5I�"9�؝����[��`m7��î�WL-�6��>�^��!�:]�{�W����jI=����O�T��$��(^Ӧ�֎l��l��Y��
�S���5.&k�9��eF��(�?r�A�� ,��_viS�K�8n�S��6���e���*�<��(�.`����,$�U��0[��G⒉� &�r�ŐQ�#\�2���:B��W�r<��gT���fQ��p�؅چ�2K#�_<�M�,I�x���Hi�`�t�HŘt&�WD���H�}�o��Fm��S ������_68���\TܷX�|��z��Y�r>H��9��wu�NP���0>��DC;L�0H^yި����e��>��dqq^�"�Y�]����?
��� .���I".e�ܗoM:�Ϋ_@Ȱ��-{�h�1�2�Ji���F�aʾfm*l���w�{F�1��v�u੏�YЫ�Z�c���<1^���i��kZ��O��Ҥ:��񟄡�:iba�����</Ob�,��p��NY7(���n-�0xT't-�
�h�����X����!�֪$����!l�/�|J�_�C#(�;�A-�X���ب�5�뜮�2�	y�8\/��&�Dg'm+VpF�%�����z���R"�iC�3E4��k�Ey��W�&K�y�����q� TfKYGx�d��:.�������6G���>�"��ރ"�}s�k�f4�,	b�q�ؒ�b3w�ixl�Yx��b7f2r��r�.�:�«84�3-C�����#�rX\��qܱ�8"�r�!/���Ls��V*|���v��u�.�0��w<��*ybO5�lo���{�`�Q ^& K|�G�։U����l����(kA�S�m��l@:#J7Uxgt�N��9�xM�L�}�쌡:���ap��z�S���i��b�(˶C��������4�t3�-4{�)4ϭգ���Z(V�IB�t�&y��ʠ%OΤ/��5�)��2 ����M�gX��hҘ<c
�������?y3%vᏴ��g�����������x��
s��*oX`E1O��SlĴ]O�xH�0�{:24}���xV�֢�`q���*vz��yƞ6X>f�3�M�$�w�)&=1�Ɵ���C�v������c�3�E 8|�ø��&�K�%�`���L��J��M���k-2��P�3�u��m\�lv�v�d�Q��?cX>܎q}��\�C�ŸɄa�w����Bb�V@@ui��E�;[XA1�v�"��`�ӷ��y�)��|X�z}.̔8��<z�*}�/D�d�b1����t\�\�<QA5�Z>�_`ݩ�U��ݩ�5k���._*>3���as�.��U�[	�x:f�׶�>$�4�M�+�e|g"g�_����1d�-s?�(�(�e�ʏW�E�)9����d=[ ���F���ZU�ЋϓrI%1
�W�f�7	���}8���n�0��;���tQ��Cz�tm����-~���W؜��7V����y;^s{R����S�P]?c3��Ç͛NYŶ�Pg4��0+71��,��3
a�,�O&��@ampSl�����"{58E[d�`�ٺ�w�� �d�\�_��X�O�OJ��{f�?��p8k;+�Q-Ji%i'�� 07�w:�꫎���HEc��3L�rT���2FW���W=2l�}�&�P�[n�Dfj=��=�o�@�H;�&�u,첢w�o
Gl�i�Kۢ�̓F�P!�O%�P?Z�dh6���;�ݱT��$�&���d\�+]ﰔ�ٽ�حfȧ��85-�4Iw*�I�AZ�Θ�*�ς6&��62���,��ѣk([�DNv����CSWL�p>�= ��vʾ.�
s�:��zڞG:����i-A2}Uu���t4��{�ot�B�ٶ9o/��F�%� ����{�ӂ��$�J��0Y�k�&W�ٹ�{��Y3����8}�Xނz�x�����6[��o&�U�J��tW���KM������D_T�9z���������;_4b���}U�Y�F:���f�&��ɘV�QZE���`ύq;�
��.R6�6�}@��n8�X&V�Znbqyy< �1�GH��4W8r�O[p�@�9�ޱ�L��O�A����),s��k_���/#p8ػ�.C �Z���R?ݞI,��b��cZ;:��N��u���V��:����Jה���ۼ'�u)�E�+��L�@��[�$�8�¥i�s<c~@ �
p�t�>��w>	R�K�V񲩎��� S�:�'���G����6o��$��K.0!�Դ����3�w",`b�`�yl����H5܍#����gm�Wq��0�-sż]�D�]n ��Z{ƌ�չ���2��Dr��oo	sb�S�{�, ��E��� U��7G���E\҅ͥ�C7��Cj��ZjvD���"�C�`��>EH`,Ԋ��4@\��C�� �	�z�]�tG{��&6�6l�0�M�zNlU!��(�\-�|d���f����(������#��w}�P���ΚD�M;�w�a�0�y�*��E���^�t���\i݀Q&O�7i9
�������X�0�v��G�͸�Ƿ��\����{l1ĒK~AW��1%_���A,)����X�L��=�I��B�'�-g�c|n-���Ve���@�5-b�g�w�A��P�2�5��m[�����'�u�S=�݄2�]\�'�E���̮-v��'�3R��i}��J�B=l�H���ǈ7+V��㣟>���'H7 �5	�������]�Vg)U� e�A�Ѹ���A�̘YER	�6��^.�c�Pѭ������ӷ ������HjXw� ��^�	�M���g�����IS�����]ޓX�r#| |�nt���<t;:Z��=Iew�+'Ʉ��Hf��)K u� �\_<�'��BZ�+�/!V��M��h2���a��%�I�,��U�= ��YN��P��Wi�e� _p�=����9�]�R����.h,4���~��Q�X��Ťz��B����}10�m�KD�=��Z��dHHu��H[���\6���6.�՛⾉�r�61��72UItLh�%�y�H��I�fπ���/�-�Ӣ�K�&�ܥ&���rU���{���U-��Q�>�p��.~��,��8G�B�2���h�zyä��
���^X��/Ⱦ�g�3"ן�Zϊ!�Z?Q�
>�.z[����эa�������ߚ����(�̒�ې�A:M"��he���EUD��/N#�z�$t��,{D�,�=.��t�hRX0���s�hĺ�=�p����U�i�5�=�(T�vu����cD�ׂ{{�����Ma}��=��!�Ǭ�5y-Cy���%]���
��OaE���4�}��p8́�P��d�3����\ʺ=� ���Q�s�N�A�7MF�3��f�E�Hf�x�nO\��-��u�!��?� \O����c*�X,<��	�s�"<Ԝ�F�I������T5Φ��'�\H��1X`�L�GǕ}[���.�j��=��n����:��e�f�#�V�,�����G�.j��\����3�<��?�,��ĔL��CP8R����C�7�ǔ���Q	-�~�7�nl��SՖ��\篟��T Qᩜkh�jkTn�n�F�6��J�:�$ROS{`�����@����'.�z��۞ǹ_�v�D`a��q0��%�qq���룳�����Eȅ�/`�T.�I�7��=or
� 1�Z�kmh�`���_�*��.�
@��i�&�{;^
K2k�96&�^K'쉁����^�v�@D&�"�iV�Z�� P��F��Ti3��]�h�W$)��'�HtU[� D�y��#���=�3V�%t 
_ޕ�|�א�o���_=���3s�ڳf�?���5�<�.+�b���B�1}�Q�J̺�I֕]�7�͝�M4��CUޣ�R��|��
�:�!uM(��c0��껽c���Sd-���F����?lD�=�_��r����ù��y�8!�]�<���\rK�#�Es �n��B��
�8�^��7XaM�B������<��� #�<�x�ء9�o~fg�2Q"^�a�i6��Rg�\H�M��U�p�/�����ӑc�2-�xJ��8�-dˮ6Xv�W,�cY��!xI��}t?��#'r��Žw��԰�]��A:�X��t��@��]���4X$�O�j>U�D�|�[~g���ȂX�y$P�Xl���)��u|�?^{�vS�����(��٧�9�/;H���.����J���l�$Eɧ[Ky�������D�R�	�]u212P'v7���X�I/�h��e`���rܾP(�K��t,�j��8v~V����+���V2��E�~1�[�{D���f�	�P+g��y,��[��𱚽��{���(�o��f�{W��q�f�:[G���k�I�1M�# 2H�}̱�V�m !=�谡9�y>0o�-�b��)���ǲf�����[x��Do7��ad�#-�-�)�N����\�L���7�"+W���-���_"O3�KY������*qE^?��n�N��`��� ��rvb2�������&/��OʏlX���gP6�P�Tq߾^
��~h K���8�	� i�ˬEZ폂!�	�e�*����nK�(�:�V}zs�&gq�+�J��y2��� 9�̙��XWy
^^1�&��3*J�$ V�NN��HMQH�?�!T��+V
��}��UIH�+��?�ై��c���=��S+�Q �,j{7�l��Р���0h�5a`���H3�:�l���b�@�1�I��k�ₙ���2�iܝ�-H�E��טnm/*O�u�P%� 0�I��T)�=�w]KEs��R��4$��d\.��(H� ��7�|��o_�}B��K�л�j�2V�#��p��A��oI���B�vQr�V�χ�ʢ�Ub2AdӚ��f�ȶg���\��J�}�ړSIp~2*[F�����`�o]��<SN�Fi"}Dr?����sW��鼺�����=Ը{���8бc�=Z�0nn�}�ܩ����6��b��?�Ǵ��Eo�1�¹Uɀ9���]Ĥ��P�	h��.a��=y�S�M�=W���_��U�b��6��N���Y�a:�O�OuM���2}u��!L5�E�������i�Y���q#L�'���b���3(I,e��5�9�߀F8r�#(9wdm�QW����k�s�MY�1���3b9AΗ���r�,% ��v砏4_�,(�-��p( }PP����-z�6�,O�U(
�/�'�p ��{5����h��'��!�'8lO;��SԎ� �w��]�vH#Ԅ��L?���� E#�+�Sv��@W������n
QI �V�'�a 2F$5�1��Pm���T��(�Q�Z�����9�=����}q�ُ-Pl��r��he/��B�j>]:*2z���b�u�K-��#�I������\c�^�S��vd���X�}EGSB�9������0�.�d��d�`Vq�x�u����T䞰�ǁ��+͛_��뫕�Uk�P�8�u'��ޯ+��%S�m�rYѫ0s�4����ػ�%b�=^Y~��"�>�X"��7E1Z���W�ce�I��Zp)�r�o3n2'���U��T�C��tKw3���E-E�i-҅t��G�X��1z*F{�j9�k�	ἂ�Ⱦ��!�d����7�G��%�q�x�`
$
c|(�y���TU�=r}ˋԻ3�g8+���:�����%��aA\G�D }�k�Z��ܚ��{W�t�JqGݩM�)XZ��hA�N�Yѻ�)�
����cu���w˔K".��6��!�
aa/�DX���sBI�^BK�����w�m�o\9� �}�o;�H��F��~(OT�|�����9G؃<Q8�@���`zR���s�ȱeJUM;vR-��uwg$v�UK�$5ʱ�+!Z���3���j���ؕ��鋔}�9�|�ێƌ�����2��#m.��VY�i�j}D;�����p����<<7�{�=9e�5�&�5��2�H�`L��YLy�3���b��x�'EW�J�\}��GY��S`�&���Q;!�[I8vLĸ?6T�Dl�=���ȑ�k7|�\��Yh~�ˆ�1����:_���Ţ+�<�b���Q�g+F�_�~? ��8�aF-��Sإ��k�|wQ:��H�i=P��FGI�#6����o��=�����G���ڬ�
���-�<Ot�K�br;(v�Xf�!��l5��9��W����c�x�^�J
M�q��W�1�S��IV�e��=� ���a>�Iq�q!AS�J�啱�l��<�߶�FZk�X�/z�g���3�|HZ�dzE��mJ�����A���ҕ��`^�>	��^)O������?��8�:�L���N��G�;�'�t�|y�M����k����}����h���I��:�Ѥ\��Py럟8eS�����K�J��;�F�64d2E��_�ٶ�`YS�j|�/6�����6��t#m`Qv�j#{���g�Uh��3H�j�zԀ�e	�t2Gbf��UP��R���A�N�!m�+���������VI%��;3r�0<�����Q�(�߀ou�7pA2;����[�C���ݡ�x^��k����]���pQS)h�3�/�S��R꺅폖�q�-�<�B��0/~!��U���\�CX>��˿8�q�=�|좖Ǫ���vk��4�1��~�c�l�x���n��]-����:M� ���`��7�,�,y��#�R��;m�m�+�d�j�aC~��m�n6��n�8a��
���AŚ�W]6�Cd��b3�XKt��q�08vY�x�������[(��^����~�����c�D)��º{��Ƹ��N��"v܈�'�.�<�CA6V ������eb+�?�\�3!��u���s@�*f�qH�H9ބ�-O�T{�BG�����_b�h!�ϸ�ij}���/H��9N�e�5��V�" =/�8[e�^�(�e�m���SJDWx~XXB*V�4��An��9(�
�?�̥jaRį�W�:�}�����}��+�9��'���A��r�N�Y�A�����;"� �y���<���>g�k}HM�"RҤMްD]b�"V��,�T�{ݶ��O�gV�r�_ب»�����$�v=#�a�t'bY���kUm��B7I���^����慪�m*<O^�W�<��~�|m9�H���Z�
�}��%��Y����7����r^)S��X����3��碸����)�hC\*k[7���n�f�T��~���B�0�=}��3����م�aG��s���-�C�9��2_g(��Yj�W��M�E�1*;����A*�Q]��]�	<�� ��5��2�г�3�I���f2|��S`�*4--��[[������f�m��D�kU+���b��"��̔�͜SQ��(0z+�q����3I�`�o+g��H�u��-j�tKvazB*��M/pMˏ�*[[��+5ɇ}^��S����9���9�ۥ oJ���T�#��A��y��鸃q,R�� ��*X�z��#����?�ѷ��T�b�!U���,��;(����Atp���I�� ��`{𩲚�՚A�AA�sn�cW%�Ε�f�M����[b?d��Ԙ4ύ+H&n֐���k��1�(C���F��a�k�}��w��b��j$,z�y���� ���,���Wl:j1��S�����c��Y�DP?r/	qpF#Lb�)��LT�@o]��Dq�ל�Ff�27zO��d��Z]��;�,su��FgJ��߂��d�q���Զ���Ȏ�t7��R����yN��zݸ��gW[������� ͼn}D�&�)��r�W�Nv��O�*�x��NZ�0��R��G��b�|;�U}ĕ$>�b�i��-$��ae�R���{�u��9���]�\�X�ka=�e����ӽ��R�����ލm��gLʼO(��h#E�d'�Zq�Mi9r'�ܴ��>��E��.�ʦ���	���.>��9�8��$�7��K�P�\�O�<�e��ځ�iX$jj���"���\��~����n �թ5���l�%ו ���0�����	ߩ;]��g`/�7�H�3-��y�7�V/e�>��G�8�t�nz�Hs���Q�rI�<�N̓)0�Z�����"L�	p���&��]�p~��àm<��akT܏���P7�:�D��Z�V߈�߲��.E�{�K��U�*
�����s8�i�|	
k�Ⅻ��.��Q�O��N�l7��犴_BJ ����d��c;���Z�I$ Ta���ۅ�ps+P/�Y��pX�2y��Bx{ ����{����s��	���j��w�m��Ľ�rm� %��"��9E K��aIw��::x��&JiN��7�'�G�*Uԧ��gNȸ�ٺ������)(�1�Y]�;4&�IFH-�ւ�$�`C��x�@^f40��>}�2�ƪS5�If���'윕�M�LA����7-ЂɄ���1�rQ/�G�,ы��v��.X��H�cv�R���Su�
���@@,8����5����kZ�%���P8��sz-zr�B�~Q<�s���D�Y���P� FC$��-�%��`Z.�ǳ�������Ѣ��h��rL����i ���ߺ���a���<RX��	��S�V�Z3�KV�L�J6��8,O	�	��]}�o� LE�2"�@Ҫ��n4o&ˤs�����`�Hb�GY���5�A폄gp�����S;]q�t���d�hk:��Sf$��4�ݳ,}��e�|~�eo���g�7�{\��)�����E�ò_u�ȡͧ�-��˵��a�cPzZ�ŋ�w����]���-.�*�_)x�w�(z��؎�T+�J���/��,��j�c$s�"ۧ�T�7V�v��P�N��
d�	B38V����n}��у�(<�-򅁉��&҃~#G�GF6���F�W���_;d�O>�;"��dհ|�eܢ�?iٞ�)���A�]Ric\	�cW�{)$���u(|�x2!<�]��a�PZ��xf.�Ԏ�/��\/.?�q�U�m�g�Y�A�#�kV�������1ё�QGP��45���i����i:_`�Ɉp�_(�x�b�O�����x*�<=���v�n�Q��vm�W��E>��Q?Чi��Í�3O���<�n�̀�sE������>QuX�4K��b�?}��27s�y�f�7�/���#X�U+���պʀ�;�O\c"N��a�vt;)�z�����ಉ|���:��?�i��9;V�8l�D#݌2���n
�L<��-D��jTwdy���!�{ K&<�����&u.[X�D�7�)w�������1�j��
:N��Is�oƲ�c����Q�}$��)z l�I����q"hEއ������"��H:��?��J"�g_�isx%cn�&ǳG��g=}���?�
�~z�5HG���[y�Ca��;�NQ�S�܉hw�ww�!o��g�v"²#hq�=�B#�]V�l�x���?s~>\g�6���s����0`���J9�|�s�!��L��!����������x��#��ԞM�ٷ�NUOr���ZB�t����h�Yb^ů$ � J��ye��Hoж�����j�L�HG�������{(ծ���9(�D�]5R%��ϋ�����~����	�0(��m)S�8�E݃����I�L#���)��y�$Ԉ�DթrN$(,	"]���8E�w�>ݳ����]͸[G��$�j^�C��\��'*��H�R�(Ӏ���er�,1D��\���#�+����r�rKA�Z�;�$�9�$ޖz�34�cw�����1]7� k�����*���E�d�ZB��zh���:�$���aR��^��@��CO����7��6+R�[%�+��Ga g�E��� [�Q�Q��6P:�"�ae4�S��<�۲6On����3�<�{������/�*5'���T�9�5���s�:�|8�'�Me��H�v�\��p��*@��*C�qL���#+��h��ɷ���>n;�_�l+��1����n��P}MX�����N��0wQ<��*1)��E8�b�(�B� �T��H��z�ԊL��˶���u��ko,y�ȶ�DR�
N�9��4��Ƹ|�p�u^oP�fL�!/�v�ū�]?y��Z�1��C�r�C�V����HG蕚y����N��j��ʯ�a4�${!S��_{Vle����48��3Ύ�-�b�����R�5P�S�O^�vP��A�]���oK*"�?���H���^����p&�{;�ͫ+�j�L�f��M��_� �k��r���v�˷x�ui�ƍ����R�#���b�h4�{��z��	�Gg�ǈ�3L(�g-�-/���>
���DyX��?
GҹF<`�5��C.���24q����)���;`_#0���\N&����wy���GP1rT�^n�'�[lBN#
��Ϛ��7.�#<��m�_;���B�:�������0�jk�6��}�y��ؿ��;��f�4��\�mr5��+<s:7p���@���\T�i��J�8�R�!��#�Ё��=��B�����lY�n�;�^���d��&N`�KT�Κ�*�]�N�G�O��;�?����X)y,���d�TrI*���L�C\�)��e���Q7�j̈��»P�S�h��V<`3�a��X�M\��	)S`��1�*�<ɿ����d�G��[h�4C�7Du��.�T�t�xy�_� k(P�)e��pN�.��W�I	��50��x����ث@ѳ��?]M�߃�����<���HU0�� RT(��m~d��DSH��TNy���@>��!xY���g�5?m�xrZӆ���\�TW����:��I��2$�4u�BQ�t�,u׎^����	_��d���ɀ����ER
�&���;g��r0�3x�k��?�� P�ݗX������q4�$�C�uAw�W{���s屃-EǕ������3󞆐h�:�[��g�+�B1�-8G9�fp������:^���exCYb	�8ޓ�I!W̩
�����?QCV�nH'�
�Uʜ��u�t����
�'��?�$)#��I�[	�������@��G��͎�TL���_��p
�|,1�6v��C���a�ftݾ�c�J����B]Otl����Rm���9x��I_ۛA��\/[N30�C�Q��P(W�<�[����c���d�x]��Cهp �&T��S�7պ!�c= "�؍CfT��(���9����y�4�7��=�:KA�['�|�ȏ*��,�&��m�uD�
���ve��"3[3��hώ\�R�T�ڍ��뮸�0`N��}� "��u
���f7������9���w*B��Ud���K���)2%�lM�.�2�z��{��Lv�� d�1'
�M�k�*#�c&%Z;x��ǻ�����H2ۭ�qv��԰l7 ;���6��6��|&��c4D�C�����Ƹ���u����q���H���cR&uX��]������@dg=��>6V�E'�xs\��e�y��V�pl�腏��B")"������Գ;�����	��!��D
x��5���uZ\�0�Y�#�6Jm��$� #j�Jx��G��K�&�pѲ������|G�vo̻\ݙ��r؄d�C#e��\]i&���7R�o�EO�^��Q�]d��ii�Mߍ��7#}h�;�`��Rz��4���7�5�2*u[�V����,�\|���a����g��3Tip?Ui4�q���f���p^�Wm�aX8��i�Z1ϱ�P�D'�=&zۃ��
��m}��PnKܰe"����k� �\_|0�m�l�N�Lf�f�C�L`lV$�H2�����e��Ȁ�����q�m%s0�/m���[ϲB�v�Q�Q�Bv b���PP9�9�����õG@��\���K2#�o{�i^��^��b�sd��lu;��dL�����n�ϥ���c�͇'S��P��P��D2͗�br���y[��(�Bq���w�a��dʅ�=�\i���́�J�X�&���:��v���eQS����:䤰z�6�$��o�ؐP6��9;�M�����)G�U�;���t:m3`@��P��9i!g������7�L\��(��]��2�a�#���A*���h.���eK��t�*Z�?���ʜ��[6�
&Ե}��:
"(3��TA�K|XF�����E�Z���%��l4���ձE���� F�JX�K9֬� 
�����s����]��:�j���r�����i�k)�1zY���ƍvU^,��]E�F6A�w''M_�F*���>��|>�1�œ�
���@@㴨,��Mh�)u� $4��|�v�����:'�-խ&��on�hՎJG��U%	:0K;q-/Z�bmʍ��-<�Hq��$����S�I�ő5��e��R�Gsˣa+|�6��2�9���ٯL�4�w�{)�	?�S�8���7�$9��
��m+J)���/��()�UV�;�zG20 GT�W��X�6��	&�+څ�$6�v
[O��-= v�G�9���wΣe�$���42��o��a��=�DD���{=���x�2��S�2���A��v�~�6Wg�"��	��b~J�>�0[�T3k�TV�>��vw�Y*�e����?!�	������IN�P��9+L���]�%�P���+�
����^r�R�8��}��0��XOB�h]�����Z��pL�c�H���W���N�R'u�&��t-��3Ӻ�C�6��D�e�D0���$��]�u�?�TS����p���M��B�^��
=N��⽄�(�$�gw=_(��y��X��W�Y��j�q2��H_���cR�ĝ�7��G��D¼�[)m|�T~,�9_���g�+nN�>�/�Χ�r������}�8�fs�u}���@{;��?i����"�l�tr!�d�mG�����W�4��_U8��yナ�1�!>���o�R����� W�*w?�*Ƃ�Zem�#`�J�'�U�ǅ���7�d�s4�l����{a�D�}1Bŝ����u�R�%����7*�B�=D��v�Yj�[�ڵK�qM-4����G�[@�'/�Pm�Sj��V����*�=�8���q��[�~�X�U�Xm�FV�K�;+�� �p���]P|�7[�}|x�R	�!d�O���d`jՂƂ׀��^�
��6$sMG�7ʾ��Q����TP��
�蚻Zp\�狜�U[y8/�lJ�}d�:�2�%j�]pj��uw��5L�?��Ȟ�ǽv����pUg4^Wl�u������)��Æ�Fz�[f:/�V*��_�GUm��h��k�9�b8��m�qy$�	��-[�D�o ��8�?��G��� m��[iC^?&F��~���.4!'��h�C�&RY߱qp��d:7p�r�+��̤���;V�껕5/�Z=�͜N,^<�����/������Ƭ�h���t|�!�6(�AУ�ōG�E0J��xv�
tA��ODEe��� ��̡��&[��I���SIσ>y�>�K�rp�������Έ���#p�ĥ�L���9�"p���zX�"g���0n�u)�d��ـ�c�)2䤚9pnO�gأ��|m鶋��4��Ӫ
��[>$����@�! �j�qz١����P)U��yk�рFX��]���ܮ�p4��0������ll���W�.�QO����aV�eG,S��C�³7����vb,S�Obٶ�E5��H�l� m���-"pJ�!r�8A�qF�b��6��2��W����fItl0�F�2�	[Ђq�=�,���\�A#;͈j��=�ԁȳ��1>2D��POp�oE+Z_^��MCHV=Lrk�a�d�)-CFz�EEi�B�$ޛɎ^9{�鈘�ܫ0�m��Q[�����%�'�u���I����]�╚���D�3*�l�E�Q<��gL��@��X`j2���S*&��6:ծ�.{{Oc�V
0Ů�U'"�b6A�Qx�i��漮>(K����m3��m��Obtg�+!]ʛ�^ܜ;��u��3��f �vH<V��m�F���5�����mR��"�J�@P��Q��-�(_*NS�lMgY�V3ny�5+#�o�!B;�yU�,� 
�>9HS�9ˍB�"v,�l�π�Y>K���5���=�
 �����W~x�2��+W'$z\�~F�K�p��������(ڶ��}�I$gd�@�!":C}L��-��<�R�@��_�7yo9aAQ+h�,��ُ<�$
4�{B%��}W�ڏ���Q5Cjɻ@(�T=���}��je�Xc2�yR��څ��i��vZ@y+���x^�hjᵐ����X�@h�m�Ahu=g+p��"0(7c��	A�ߡ2�ДC�N�t1:���k�N���K��J�������gy��e��s����.�l��eF�3� �&:����_���y�'+g$�XM��$���p�i�~�YO���<a
4��>h���s�e�0)��}��("�w!�� ^�x�DIM����{u�	;���k���tq؏�8`��g���/�ړ�e";��]�Y�Ł-U�*hE%�)֐��@e��d<�}��n�С�CUv�ɭ~������>r��-��α���73���| c;?��E�"����]� G>��fs!(��(7ZE'Kyвh����]�a�.�ɫx~�B_�(c��x�rk�n����2{��5�T�����SY��?�G/s�e
�Z��vX�$ˠ�\u�S�j'���*T;	e�P�s���)</� -����2s�R��\��N�K�-�gG�~jvx�}Vr
�/$4�Q?�~���I�ݻ��B2�!��F���q���-q��l��ǽ�����N�1C\>(�̞j�D����ҿ�g��,]TC�]uaȁ֓4u���{qԡ:�1U`?�An��T���}>'��;�4����Y+zz�t�v���ց5_��$���t���B9-A�wC�U$[����J��?	�z�?x5$�܍��z�#Ar��w&�o����{��,��Ib�j,bKDw�rܛL6�<*�L�ɞʟ� d,#ױ������u���pb��|w��z����|��3���k-K�x�9V���o#��~Sk� ��}w���m[h�r�%Iy=�n�W�P~ʣ,x#�V�>i��ry����e<�����H QƜ곁�8�¿>���R���� �� }�n6r<�򡒉�`
�o�����a�	֗�j�����G(��m0h7s�y�����o���i�m�dh�G�F�������>�\)t<�m���4e�=`4��"�Nq�3�^�=o�T0�d��e�b�6m<uu��9�ơ}�t�LOX�ܫ�a�"�+b����\r�|������ǡ�1p��q6�37Z"-��5��m!�h�mˈ�V9~�y�G�2��"�Y5��3Fy�}�c�n�tPÙQ|��]��=�n$���0��1���y*�;���E���n�K�Է������Td}C�G٫����fƼ������(���31��"����Zi�C�LS�%�^�O���<�l��K���jh��ӄ@qNO��F<�����<ڹ��''���O�C��Sr
n+W���O9�'��$��@�]72����*�e�]����/���F^v7s�n}���iYʝ�#�F�b�w8�{��kp6�@�͜��7CZ�O�T�G]u'��ڒ)�S�@ުy3_lK_'{�Ȑ΀'�>@@r;8Kb�4�
6,e;�V�&R)Z���^��E.���%���h;	(qT��!,��z˺�I"�f�<���kH��aU"�9����o ���F-���ʗ���{�Պ��'W��Ϯ�S�5��
������f	��ʺ��ċ��(R�+�_d����r��g���(�ý��h�C�ܯ� �=>�S\��t<٫����Qr+Vk�fH.?]{i�8����^�Z^�m@k�_=��̤d@�p�{��:���*����nԈ�.��@ʠan��z�~�z@��Mt��O������7��P��欐c>�쏋;y��NTc�Q��R�����Xj�Y���J�-]��"�r�Km���v`q|����v�pdC������
7�<{!���eZ���ks��ߡ�U:? ����^ �^#hь�i���hk��dT8GD��9'A]v�ʯ���@.ru[�'���ks��/Q���v+ԡ>�(9��4N�	ˇz��"�����/���5����?,n���Q�<L@���ȿ����,Q��2� �'�hf��]��N�I�ԏ��:�!}�Gz�◍^C�N�Y����`�@(�{�bi�UNv���3���;5�o��h�[�������=��BK#��#i������'�Ђ�?v5��A�QuzTI���V�Dw!�NJE+_��^,�e<�v��1��L��遨c�5�a툵��O�?=�n\��F�v�Y��h@��}��VE�v121����@`Z�
%D��'a#U�V�M��άɔϖ��!�@��G��5x�4��(d8C�JiX�Pn?� 0i�/޳P& �E-?��^7�M�L(�(���"&+����!͒��;�w+a�2��x0�߰��=]2&^y:}ޢ��qA5x��R������C*-��C�oJ������T9<��v�o�MK�HL-uyJ|&�(����26��K��T���ԗ��uۋ�7�t���w�Zg�q���й
L�,�R�������*�p71�����m%��}XE`.<iAߧ�2�j��)s�2�$�!�梯��#K-�K��Y91�7�*|i�H|�a��@������[�vu96�́��Y��� ��e�~�i��[��!��kGV��*�����J
�i��eq.����u���F��dϝ��������p���~L�]D1𥒽�F=)�|�;A
�HRT��W��^�Dmk��3�5�8���ūa�����h�ω7�wb,�6�*(k}�_׺����9J��<��:����ޱYێfD�|)�y��L��!����i�)xz��l�e�Reo�ѷY:�_j �ڌ(e��̈�4aQ/�H��S�����Q�z�����@i����?D�\}$9������)r�܉&ل����(��Y��+��w�/��" �lIbZ�9�hwﻊ�_ �&�?,v ������Ol(g��ؔ`N
��&��	��s������}���M���XP��V�q�R5k�ۑ��w9T	ÈIݿ!HTt�M:���(�I���̷f\���&x�uE_�J�'L�ؼ�����i9��ԣx>���� �I��e;u�R/�7O<���ԯ��1*d9��N/Cr̽�!�8��]u��6�F������o�������u���$�=P�Ž.�p��b��_([��"[�:��6S*eI,_ODF��#@#-���\�/��"��
���h��+�cr <ڥ�MȲ0F9I�E.��]:r}��T�_	��ѹG�F��ի��T�a������ȷO>XB�������ܖ�ɀ��.-��㧨'e���������ELJĄ�^!�f��˿\ۻH[�9��i4�'~�|`�����9�i��t�S����c����qq���d?\���_o}���O ^(�˕ͣ�Xd!?��*X	��������/6cA��,?G��4h)(G-!�2G�Y52q�q�aϻ�yC����
�����$�$7W�R/�$�j�~J�n:�J���I�'%U����(.;9[^*�,N|u�����0����[�	�#���W��[�[����/������&2��um�h����}H���&��ǘp�Pu�ҷ����ҳ8�ϼ2q�����>[Fa��j�8Y)��Cj�(�h�j;b�f���o�a�AD�dt����L�W`I�s���d�N�~93���Dz�j��H�Z�$7�N$w^K(z�eDi-��}��q.�7���v9ϴc��G	�ЕE��|�p'%{Ś���@��m�:e��KL��NWL��Ԅ�����Q�'kF�O^{?�8'��R���6C��ڜ׬dL��J�y��qnk�a�L�M���b;�%Q������T�?,0����aao�L�����QS���ɛ?��N4�ׇƎ��d��E�ݾ�.Y9�w?l�͋7e�!=@�o0�LmU��k�ӆ�y���i�R���m�phM���%9\�:��b)���A��M�� ����m	�u��a��BJkN�7�j��\�����9�O1��*���=>�XL�[�AnpO�H!���7 p:��P�Y�z��y���+O�r�����ke"�Vncm�r
�KK�éB�vN{}��6�T�����N=��HP}\`�9��I�߬Q��"V��-[7WPx$��x�����
�L3��`$�v�����#%��Qy;���N�6���_|,�O�%2��*��$d�����t?���C�IE70L�eI���	��r�A��V��@�g.|9�K h��3iK�Ea���"g ɟ�t�\�l��� D'y
	�A��9��zϥ2�$ܻ@��0���9������00>�G�4Z�����$��᧘KDI������8�N*W��'hJ��%,!��q�9�A�q�z����9��5�8���E��­��4�;z�΅��K,�w�R�-o�S=��@�LC�S�R5�����B��̷�P��6�^�WE(i0�.�S�lF޽s�9���d�$�ܑ~p	��|H`yW�$�;T|q�y
��	��y��������\;�.--RZ�n�¦b�C��f*������o�k����Ω�;����
L���n��6�$j3�?���<���Q�D��U:;�BU	���s�0��r�:lw=T�����H|����c�Lr-�s� �x4}���&��	X{4h'�q�����D��u�ro�>G�{�K�7��~��E�P|y��f� Pt�X^!R�#�I�֒��W�X��,��(�	K��5EX��,�+�Z�z�+��$�8���K1����gY�U�'3P�@A�T-���L(����)?�ƺ�h.�v��S���}����r$���$��K)N��p�c���lWz9Yz N��i�����!�]M0�ڈ�\xob�%)�q{�!���P�d�D��;���?�O�{�AH��"��8�K!5+���⮞;�{�%ҩq����B`.(��߆�s��9{��F��f8���j@F��*���R���5*���,<w��}���<I�!�
-t�b�$����$c�HQ��'�����}��A�le�i�nӀ��!M��b׿pc[��9���O���^���+vc�%�Z}����2G�3����ƉFi�+;2['�^�U�^���5�]��l�O��̲�7Er�Q�#�p�>k_���-��=� JU��\
ok4�48H�� �6�4�z�J�TP:���VK��?�)4�24�5��d���U0�tV�
���R��3���O	O5o͜�����z�v��c�|pfDY�{�}������:R��/������F����Z��"R0�BJ�9����1��U���V| W~a�(s���T�K���W��7���+[�W�Ì�����kv��Mʰ�"�(~�k�?B��g��P5D+Pl3�ER+�Z��%� � qQ:��ᬮ$�ڂb)G:���2�NgRD�"N��{�N��N�51���X6NOԴӒC�ؐ�����t��A@z�M��z�Z�SY	�TK<l&x�(F#!�9��c�����jp<��g�2#�IP��D5#��z\1L:�U�g���ʙ���p,��}?������k��Hv�`�A��:��$�)= ?����SSd�Jw�3�)\F�j��DI�+�r2��5�=֟��e�i�=�Zbѻ���;b7�*�?�k�~~��_R6��[@0NH�W
���X8�Ŋ�\��u����&��C6��#xm����j�z�����ݙ���
Nb��.�O� �_�2�?Jas�ߔ5={��qzq�v�`�s��=�S�8Q�ӏL��Ul�R��n"�
Һe��Bn���r��=��g�#/4؈�9���"bi�@�*6vAe�c?Iv�Z����K����̓r�o���w�|�AC(�r�������$í�����ee��[R�Z^�+��l�7m���W�N�T�ud'A|�}�?��Gl�g�`[�_���s�n�lW���3�����ᯒ/(ү�Hd�B����J\D��|C:vS�:t�5�Q��y�'��#��6C��[.\;g{���+[nt�����ū=l� �<�J�`ޜgl�)���MN��zU^�uF%��]���L�~�xT#�z�(��xE���qE��D�j%G��*ru�D�>F�&P�~yT0�;���UAw�:�Qj8�}��i��k�Bn���[,W����ᗽ��]~F��~�iX�u^��7r�������{[�}����|`DH6�Ϥk�`��k(M�II����fW� ��q��[ن�-��FH�\�!��x���#�m����L�Z�-��f絈QLS�1�8��@a�AEJ�YV��vb��
��p���.�"IP���'f|r�6�>��x�rsz=Gݹ���lӜ!�R5��p��ܫ�H�#���c&$�gL��S�,�am�>A�D�7��?��-">9'�#* ��Ah�K4ѿ
;�/����:7+��³Б~�"L�CRy[�Pc]z0�qEDê�۴5�~v�f�o��s�Tn,$e:gVV����gR˚ms��l��� .�Җ�l��2�GX"#ߤlF��p�r%Ђ�v�V<p�P|���i>��K4O��2b/������q�PeΖ�iKj�2oP݉��'���N�N���������=����ve��_�Xs�"�e[W�q�|�䍙��۵��af]з^Fk���$�{�Lj,��M�D,��b8
��m�>=D��V�)[t����*����BƏq�X9���n�DW�/{�.�3��:1�����t��F�.o*�R8�1��\�yO[3p�Eh��'e��}b%���nj��6�+��X'�};�㼺���ʊqG,��� �V۱�Nb/PՐ��tb,ͅ��Ky\���5P0ڄE>*������b�����M��Y�G������$;���L��aF��e��<��y)��߶<�Y�(=�=��ac�B������ ��ԓL�ld�3#mҤ��WR�P�1uxC�ө�mN}�MT})�GV��}�rF����q
D�R�\��8}�!�����e�ٮ�#Pڏm�����m�[!��h��/�m��e,�s�������P��h��*���t��Lݢ=6���r��A�/�{>9�|�3p��ӽ:�v��)���%v+`'���鷊�F�g ܿQ�ʨ���.d(�ȉ\+*�%#!�����TVoUP;.�����S@	��=�������Q�cٜxA^MC�#-F\�����:�jà���[����,��
M�b���wލ'�uan�+�GFM빉�dAM���?��n{y�:S͞R�*H�|�md}���3��;y��X>��i;h^�X	v��9],���_��-5�������฀0�������^2��%�=0j<���k+0�q�]�/L�LM����}|��w�B��\��&E��6���P��C����R�4�3y�.o����
W���͂�%R��[p�x�b��ٌU'�,��~"F��]����w^`O�����}羜�p1�9S�u�5љ��]"`�~��/o�$s�"�FaɄ�Ǆ��n$
���B���8l/<� ���^����.wع[�����O�q��Q�G����}���2�ƅ��S�B7��൮�](�b �T*\��LY�+|���ڡ_��������2JZ�_/�S2�W��^o�q�҃\S΂j{A���ו�K�Sr�����g��<���%�O,{����j3�u!�Ve:�c��^�6������5m 2���۝E��CgKS�}�P�x�i �rc"�z�&d�C��o� .m4��Ӝ�N�e��(w�q/�	$��?�-�e�Jk[�N�ǆ��iR88:K�8��?=� '�	#������x�.��3$=���{�g!������]���4�Q��2=�-np��Շl����H2���5gRG�@&)Zֲ�K���[���%��G�%�����Dq��Hv&t����W�H93DE�@���3O� �0��Ӽ�$�J'ĄnC;{�%���q`,�A����B��c�2��";D�U�E_B����[~ZKƯ��@�2�0m�˵��O}����:����[*խ����yV=N�A��
��w|�}�I��S��vK��;�EKt�w8#DB�f�NgN�����S�����/��"ѩ5o2X�<,�FEۍ|��cP�Ð�ZmF��ôb��b`?֬�;�F�հu�]�Y2���ݡ=��)5 ��"P?�$^�^5�����&��c��>��)w�ut�֕k�q''���:gh�9�X�O���Ɇg4�Nֆ ��x
�F����	���y��n��>���?��1U��X�qC�c�Ԕ������h0u�;S>nE�hs"%dx���9t����4(D����q�0�aZ)wa�33��b��]M��{r���"4�T���ݎ�����"��y$����8�]v/ޑ���0���~;�e<����}��c�=����wP'-�F&o��2`�`7LAHí\����J;s���Q�>���hU��B�o\�w[�Q�k���(�gx��<�s���`�%���<g���by��ǽ(�o7���<�����_^����c(�a4E�[��^:ƚ�h<���4��{��5/��[7������+��q��"���������T8�=�\�c�u�TUvg�Ml �LGj	��׽v@β���(�%���Pq�-W� Zf��%
��1��]!T��ď��A�_U�*X� ���Ժgm�$�"�U0ké&+Fz�pY����� 	t$%T�g۸�Y�#l�����>����_���'��k?2p��>��PD�~�:����B�DGt����[bݢ��1K0�` �f��n��X�s�çm�8��|*�Y��#ck.�!(����maȡ�ؠ�P�j��Q���X&w�i�PB��g+�D��Ͱ+kl�H�2#�4{�U���[����I1�+��jUdy��F��9[��$�D�/��>g�XR�����ܮ�`�! ��N�K�%��RtL>�{�P��Q���8�����ǁmδ~*|B�=�0����D�ڼ����;�҆�%]�����������q�6�d0��.w'����l�,u�50zu'�ᐎ=�-rRΈ��u}x�$�c�̙*7�S#F��P�������J�玸K�YR�Zy^�1�pWB��e�a���f�eCOg/�.(�V�Q�ԓ�U�O��Q|�A�����眩�~8J9��T�� N,n�4��J�Ϊ��"2oػ��월��9�F���������g��6M�S9�������k>rɇp��Y������	RZ��G���"�(�@b�l�+F��qrv6��|q~*4oR#&J�}�%�'���c��w`	"�슀�<�Y1���aK2��+��@�]��#���ϻ��1;�2_�K���r^ط�;��'Ma���y�)��:FSR�8~5�kܣ�
˖:�Q���lz�c�'����,��K���p��2w/.z�������_{��hz����[�4�R)��o	08��@ք\�,�,��6 �(&T)�#�wZ�fVn� �1�»R����������<�D�ш0K�X��2Y~�ktHC=��N�3�8l�����l�R(�L��F޾ ��6�x$;Q|r>�@ĵ��l/m��aC�O�������1�U�EZ�'����ް�v�����%�V-K�t�t�[�1߮�؈d
����}#����]=�乬���I�i�k�JS��bpr�*Tl�3�͹� $HZ��-M]\����AL��-�^j������7]��SUQ���&��r�©�a�1+%�X>��&��B&R�uO�t��ϔ�t(���Oq��	8��mr�'1Rz�P,#��?���:3eJ7}�C4�%] ;_Q:���Ġг/�o���������E�<�f2������e`�@a��w\�:+D�Pm���F��n�_ę���HFƍ�<B}���k2��G��ȟ��D����̍?��ZSj��-�R��0.'xu�9|sܼ�3n�.s�	�u�ԩ����V2z��}Y#�"ꬲ��6�GL���N=r \����W��ڷ������jq���%��-��Q/}���P��$;��<_j0K��g�ڵ��q�*ܝ؟��agT�h�I	C-<�X'lv,h�)��} �}T�'~�-e�y��_v��l��#	;���J��{�0�?�C�H[�ǣ���
&Y���\ֲ�z�U��>�KlX6qx�qԝ�!S�x��k�@J7�+S�Ȼ�d���"ÞF��vﮙ�ӌ��R�"��[��2~�<u_�9��=9���w��lͶ��1q`i�I��@�ٌ	��o٪��uox�0�2��ʞv��2�R�t�e��,�	�:D`j�C�&Ç����I#*W�ʶ*�dI(F��x��v��u�:��Ԍ�� �:���S�*�`T����:jQu�-��t�R���tKm5��`몋_�����?�����8	 �tv�R|<�1pV.@Տ����Wk���4ڵ��EZ�Ye�+��
җ9���"6��Q}���2����:T��j�Zy&g�%����be�G��XpX#�L j�|C���ɜa%�+���P)x̡���ԛy�n�{cr9�����ƀ�rn;�cf�VZ�"N�ǟ���Bf�Yu/���E�
w!C�
�1�����6�:�?�E�Sh�o�8�Nӎ�z:hH�¥�v�����\罙��8Tf���+�|���0OCD-��	=3���lޚ��8�QӾ����j�A��Sb�2�9,�I�����JR��8�	�`�Q��1�<UZ2���R�]���+X���*�"�("��qA��W�B鶪��V��	��nB�ϕ�k%�o�Я�(�8(�Ǡ@��w�_�\h]���B��g�܊�l/���(R$�?�qC	;���J�'R��ز~������� 4�g���AiPwcK�_�>�H�t��N�t�Qz��փ�TD}��B�yrTSD���h!����@UPf�t�7V>�9QcF+���\��eՔ�`x�C�B�O���hz��i���@r�f���5�E�A���.���u�1G�"�y ?H*�:=��''��Q�/S�n;X�����Y��y�^�0L{RFe�'��]��m��:c����V�+go��M�jWJe*f��D�t!=��%�^C��>%^�*�P�T�X4r�S/���tF�T����w�CE�|�� 3�]2��t����Mk�3Y���O��O`ؠ�������1�w�A��%�=o�K�׊���<�d�m��ʪ�>:%�[���a}p�m#���̢Uw�O�`۩2�t����gc���U:�l5,@���\����O����LN��~Kϣ< ���a���e,�D�n!�
hʹ^��x7��!�e�T	 ��YcI|ڿ[��3z��Ǌj?U��G"t�/a��EPK�}!���U�Pb7��s�;
Lh`:Le?ڍ�����H��ߏM�/T�\z t:��G|)���TdF<J���+�rWJ^F�� Q*Z9b���Mu�q�r�=�]�MU��^�R�AfH{���_	�/���/��D�^�axק�q�K�Ba������ �&aX�T(�����Z�Ѫ��5`�Ϸ�l��fJ���O�~��+W���	�Y޸ zrz�K�i���ZB����?p��yɨ�$f��/'�`a�Q"�����+�ߏB����3����gv����� �����+��f�9f����eG�/�i1ܑ�.����A��]u�eiD��N��th�Fc6��b�B��8P#��'�]O��^K!%_�z/Q �
p�6y�z)B�`-z���4φD`N�f��h�r2����:�l|W�B�������������ı���ʛ���RQ\����DQu�y��R	�f��O��M&�9@&=M̀;��e����ɅB�tC�ӕ44���ƛ�r����ԯ�)C	�Y��2!=ʋ�B,0�����!�5.�s��$���F�wZO�����s߅_v���?V��}�'�	�H�@1�SI�S���*�U��݊�-�i��j�A�[&K�::$�O �������Q_��c��Jm+B̠-D�A��9r����p�D��$(��%��.)�Z���ơK�9�Ԣ~���/�GP/��O��������/$�";�����=����y,���:��w�Tv�h�����Яش0�ƞ��^*���z*7��M�ͩ���q��t���ߩ�.�>+���(KL<���`�ϟ[t��^~bZ��X����Q+��\�����cΕKS�u;�u!zH�"q��40w���/	HU��ٱ��y�h�|������ �����Sʷ��� !�OKJ�ҨW �����P5�&��[.�x9:M��~�$�W�}��]O�����;����Fe��2)z?�]�CK�in�Q���(J�J��J����=y����+6�Э�ёг�dB;Q�t@PW�:���a/��H C�*��m�Y���wG��4���A9�VEW�r��!b>{���4S˧Ų�#F�G������-z�D�	��e����y�}:�Un�b�M�w.	�r�&M���Pjk��6��ʤ������D{�T�f{k���Rk9����o��I���D����ib��9�m��M�iw}�ؿ���ЍB JL��Y�E�o�k�Mz��d~���D��D�⒔wxy�~�f��U���C��k"c��n�����K/��E%�;���H���4��p�s=�|�:�0��$�vU9��OJ���<���8�Q�4_��۽�[,u�̽���E���\5��^02�ˀ-J+���'	�_�V�D�*Қ$2�.�S�67�!Ʀf�@�˭��9[S�<����w����rC�N��luq� �{Ώ-ٜmh%U�=�A7J�
Հ	�)�2=�ذ��0�D��u9�4���Z��"��ج���]/+�^>R$��hw~e�@x!��2"57�v��%�Ѝ&�������f�����9E@��8d����wѭ���aˬO�ZS�7HR�˻9��{�ŝ�R���%IX������/��E��Z�?���,����T��|%c����9<`rf��pt��0ݎ�H�ٓ�V�M��H�N��7�,Ї	|c�O�Ė���לK7i����z�.����U����k+�jU�)GB�B��B}Ya��c�a��$\�3q�������X4 c�� n�3��Pz{��T��e+WU;���Swk�i�;��J�h����V�+����$��;�S��G(G���y���p<�����/�鳺Ta�۽^���@�˟�в��D�0.��:uY�X�.ʅ���$W��(�W�v�>��iC�v j���&]Mf9����1��q;�2}8a������s�յd��8gg����ǆ��7fh�(-�Vr��.UA1H��F����KԽ�t��\��2��
N� I?R��u�r�� v�cF�j�6$#�p{�^#83*�+��gKhR:�˘U-%���u��wUm���$G�������5"�����ly���~�{P�Z��}%r̸8�	��0uD��6�m�k[�1���]e
N�,�ꊩ�.�����&I���S*a��Y�/���3���v@�	dG���bR��P\ǲ���$}GP���M���B�C<�����2cɩ �x� O�����Jd��,[N^.2.�4��,����oS��/����l�>f�້�{
�p����3jr��y�K&��[5�e��[���
v��g�Z/�6�XIi�/�3����2�����y�V8����bq�C�Q�?�ݻX~RQ��gn[��-eIy9�+)�1Z�{)l^L�*u�Ѐ\3�[6��k�=9�U�7��xl�^^l�P���M��1*d/���e0�����KKө:yF����O�2u�$Gyx�o� /�ʡƢU3��q�]e��*�!j���&�B��}�h�B�jAt֢�|�t�#9C��|F���l5��(�@��\��X�.�,�~ �H�D���f
A} �XO�d�,� �>T-�^mm�� ���+�0�� �L�	�\dko��3l�0�)^�3��-r�Oh�Ӫp���^�*���@%7á	��}�8�F#�RO\��~z�&E�*G�`���)d����z^������� X'M�[T8Y�<.����=���u���{"]!`���
�Y:�x�G!��w�эK�4��8�����
�� ů�0H"�5�9���K��4��4�{<�gE:�f���'u��q�k$�wffB~߯K�S�E=�S��	�,�8��mIt����m
ܧ%���m��2D]ʘit�/�p-l��%�-�b�׌��\̰}ڟ�Hk�������,�S����#�+_F���Ld� *(�m���ϒ����}���!�E
�Z�5�X��R�x����a�]^Z���T�8ڶ:vp"�Ӭ��O� >:�g_����?^Pn�!�	sF`bܿ��R���o���^��Z��EV�Q��ө(�e�4x�Pq.B�Y�\5��� ��l�a�i�)�r���{b�D�"�h�'�T����գ�����5j��h��u�~X�A��'p�-�%�m���W���dE�5�x;$_0)�_���E�z `S	�K/:��Z_x )�p̣��/ظoM.*��,��Z�6��B����
�j�X��/�%=)*��� 3�<�x-L\��1;��AC�����wx��H��߁H��%'��b�� #G�š�����x|�w[`9�C�s��"�Q{�c�n��¡�S����������fp�y��<Mn���V�&�9��"^���_��O���}���6=`�����|О��!cC�������{���_X.�� :�g�|���bp�x�g!1>��p��'E��\Ț|*�q�1E����Iy�����M|�. {wy8�D$���i쪐�9���0A�j�]p�̭�OP,2��%���Ub�� �
��=�
]\�{�����,�-B�趫�Nt}t���r��q������ �
S5;�a[�t͚I�Ģ
n�#�
�`i6��8+�8m'�x��������p� I�W���aĔAG��c^�&Mh�5.��4󂅲�Y�p����H66jW��QѴw���]�;��H�~�8�J��]����O���c0c@�,�5��m��^���9�I�R����!��/@7q��d�	֠qԥ
4��&/P������'Ɯ�-�3T+�U������|���g�ʿ�8R�%[oagƭ�>L�/`�mLwuDy>�]�E勿A��ۛ�M�Y%�#�NK��wP����s��.�����䎁JT��iȳ�#[՝�F��)�%:�W��)��rq�5g��� ����T�]�?�U�(H���B< 5��[C2����h�(���_)��Ak�$��f1���m�ŗ�m�^��i·�4Qe�3m�vl胚�B�W:�:���e���չqn,<9��1}��|�#��K+��h
qd����J����9�aEtA
--���x��K;1xtr馟
L�%~7�ر��r=��V]<
7ɩ�Vi���DGz]۹��}���-��Z+�=#	;�\BV�ؓ �8�O��{���6T?���)��%�,�@�A��� �U�zD0��N\��������{��
8�y�#��l�C6lo���\�+fl"�!brn����o�U��Tn0�T+��ݤ�N#<vrQE�k
E��R�:���$�Y�d�5��p�{����`DQ˶�S���{_zo2t|�p!�,��C`uh������?׫.o��(/���b)���  F���,I�ȷ�9�]�����`��2f�Y��^�S,�(jv��_�Z�<��`�J]ٿvz�苕�"�c�������:�%`:aΧ��c�D�c�酑zK"�<�p�+� �΢���֞f��lA�t]=�Z$��v�(�5��k)��G'J ��7m�;�6T�]���(�4�Y�a������]"��0?��V��}�с��q��X��^��*s1V�������r��� q7��|ok���H�}��ni�� Ge�>jB�����H��O�S����ڡ�I�a���Et8�|��Ciʡe����^Xk�b�֤�kk&��� [<��q]�5��KF5}�uҁa3j���+؋LR<�j�)�5��Oy�u��;�ט����c���Rr��d��PK}A�ڒ� c8�₯a'���$d6�S�#���̡�J��V3�	�o��j��8&�oֽ����d����.�MO�9�.�!ĈΫlx!��� �0F�)Э;��;yF"�x��{�W��_�X�(���-�竅2���'R�s�u�K%�躉�oU5���B�@���%)�^������y��큢С)M�K����р��&�?m�=p���\��	GW!��f����3���u�h���þ9} F���mK�7�_��(W|���g��}�Ό9���v�=�p�J�h*�@��0+8��Jљ��'��h���j�zv�D���� q�N���?700e�3�f(e��ne ;�^+�t����rR	����dR3�e��yi�չK]�������[LZ���9:w$�V�������(�0�L�s� Oe[�C�n�-�nG髆3i�G�l g��L�#���7H��ß�`s�5"��9�bv��]{rZd�;�S��.�A�(ci����T_B^wC>5����c8��M���`2TqC��]L ��w�B�p�1gaaC��.�Ja��l,��>c�Afg��#��)�]���(d��ej`q	���{�a�S������g���m$�f�c�T�u��^856|��T;;e���0}	������g�0ė���Ԯyn�ـ~��i2ϡ�R�y{z�ER� ؓ�g��ŦÑ2�'J>�^���HV5�g��{@б�.�zH��'1�3Гb��pCN1"�S뇍���p��a�&���륈��ڤ~���'��N���>J
AD�֫�h_)���`�t��Hu��h�k��6b�ɺ�V�&TI՛q��n��y�r3�r^l�@4m)�P��D����w^>+�~`Ѹ�R>��Ձ=��6<`��=Bw�����e����^�c��AY�z&�w���w�5�Y�]"؁=cKCѫ7���B�Ǩ}�/����@<R�d�D��m/΋�0h�]��qhW���A�2�,{: |}�FD�G
�ە^�n8�g*�{��wi�~�ա�#A<"1�Rx^1y��.�� �����9GP�z�8���x�E�CݯZm��S��ȱD���d�[�Q�dz8Z\��6�	뒳Zn�b�39צ�D�Rv�>�v�!�p�[�P|������ݓ�>�w���:�4n!�ya"�SNxgv�CNl��pK%�x��޽�u�F��b`��}��h{��x��PG\�W}��	�ә�K����{&��.�~&�]� rF����>��>��:̠�s�w����/�ĵ)	�J��k�2���I�ƨ����4�I���<rN8�9>��-�x���<��y(�����8ZFo�2��3a����O�G�r�x!:�q@<0=K�n^�V���S���6�ສ1�@�oc�
���vr���\A)��%e;�c�N�^�'�~����;�0<v.�����2	Rx�z��AM��ʔ�NM�q)��xޥV������ɒ��;�爷���Ϯ+j��C�3䞓��/�%[?���J(fK���4N�GSG7�C~O�F L�e3�g]Jd(�z�~ڊ&?�Ğ�OC�u�WGKq�av��1�1���/����J�3 X��P&ӹ�����Yy���^�g��ɏ[a` �p���I���{��.�{sA�DN��0��x�?:�1�x(t�UR���Eܩ��2)ȉi����2E�9@_�F�,_����#`GV�P�@�_�2��Ҫ�>�w�'0�L
�J9�~�%q����߇X��iP��ʩ�P��]%��i�l�,�O�1	zd{y�Q|����(n��f%(�GV3�N{��f6�F���!�7�Ex�9�QR?�g���+��30P�g�cq5F�l�js��#���w�:���6C,J����%�L0{�qNsk��'	h���T���;�a>� k*�*������~Ko�\��m��ϱ����8p��grR���ei �j`(z�Z�����'jO iL�PY;�Ņ/51Q�qv�w}�w-ry���'y��iѱ;�+� \�\�|yU�ye�F��Bf5�ݞ@Үt^�9Dn�O�A�)L�L���G���)�p}����Ք1�rv�布�#�T"�yc.y~ֹ�B��#���J�)������gC�/�H�T�C�)�Z|�W#<����B�� �$�V�p37!Q��	0	&M�)x���BߣF(�K����&�6'nC�qpVp4���?��"aiq���a򈭿�F�/�>0E�ū~:��0� m�C��+�З�=Qh���+�so��1-��2Ծ�zb��4����(��)�U?�~gS��qm�b���s�k9����FIE�$s)c�?�f|��I���BrE�
Q'	Mۉz��a��5J�ƽ�h�|��T:y
�[Z�� ȳ��<��f�Sܼ���-��!5��MW�L$�d<C�G0�\ȣ�9��L��ۧCWp�����.��BF��W��E�4��e�0���=�Έ��Jk��G<�AY���m�!QOX��B!�$
�mc*�G��#:cnxL�����w���'�:��R�2R��2l��4G��l��%N��ŠR���Hs�!�lg�!壥��6��"19S�</��� *y)xO�����׽A��
%X���$��C"�h�H�,	���J��|cE��.#�)��t��Ή�i�R|�V���sWg'n]!�D�V�����Z���(8��}��;��Úh��_/8֏i��<�]�-qh���?��O9/b���������L�n�j`�!�)K_�X rr��4ۨ�9�� ��W2̍p�|<�Myխ/��h30.�S0+[%d��W���7*��T/�%I_�v��W;�ϸ���i����f��Q�a cY��X����9��F��
� �+����:�p<�4Q@�.�6�9�K�]��kA �Q�_�%l�����M���{�2��S4��������_xk�p�պ�����y���RO�2�$ /���S��ej�97�}0���rsv�����L�"�^�%G�v5���E� �Gsƻ@��):H��O�Ӎh�/���̀��"�F�$��?��fr�sPB��������Y�/��+Ծ��M-C�\����V,I�0�S�X�mBS�O �{��&2^g ��K>�?|��V��PG����f��n+iY�~$c��~pgs�-�K��j�f���Sc#�	��ֵvZ �{1�\S�{]�7b�5n�!O���ziJFP�ګC��gI+b�f9,�j+/�0��	/�ˤ��k��Lr��ɽ�R{�q�\h����4���_$�x<�;��G���Nө�S�^�ǁڨt�H8*��/�V�!������}y<�߉���]�5Qm(A�� ,������c�\��;�|�ۋNe�~W��T�W�H�͖���b�Q��n"�ú��.-#�w�u\Y��NL���X��V��_7[7\�&���<?��h���f���tq��D�7(jG_����^��1��fy؀���+���$��~s+�_�q��b�X�ZN��<��>Eޅ�G�ʕ�D��,��֢�!�K�hڬCW��0��ޞX;n�_������~�s{*����@O�x���7�7r`�䉸����������P�Fe[i�B�xbf���>��|i ��;l�nH\{�H�c��嶗=���*ؠo<|+e3=�fgo���[ν��~��<��ʲ�Y�:f���p�@iOG7�={5�1Wp��>`�=�9��n]��n�����tN�vI����ܢ�u$]�z�*;		3��XM�?J/�ݮu�Eu�؉b<'��+ޑ�׋[RG���*%4�d���Y�[�d�(�(?|�:r�tRv5̱�?�E�9��������A)j����*�o!�0�Y�(���:wF�͞]~�s�R�T��\�[x堩�>�7�<m��o�J1��Z>��;xh�$�j���G��r�܊�Kx#4�1{uӁ��A	P��S�c�\��⁻l;�� 	��n>p��9�kJ���7�-(�3�	�����5�>��_tt�?� }������qA�2BaC5��(qIL���4��a�wW��4�Vjwɟ:��r��>�!W���x�����7`��W+n�G:%�߾co��Y�u�s�a�H\a�-"njL�GE��+��Qd�9[2�ݵg�~�1�����*k�Zvk�*�\�P{�'�ЉjZ�#���KW�U�(�A"Ch��/�rj���nf���m�߻M��l�݂6�sGE��lyχG�3@!vK;��e���C�B���cŴ�nj��4E,"�0�hzNn�+R����K�ŜZ�n����A�D��W9.Q������!٘b;B&{�452e@*49ߧ�'R�4�B���K�D�b�K��oR�����k�:hG��-6�!�p7��Y$��a=�Ն7G�f?̐Iǿ9�(��B��R6!=��@�B�5&���u����)w��G�"�V�Rb0�~���G�)�mu��b���g"d�n`�ހa��OR5(E���x�KXk���cZ��:]�
��WqM��(��%�E�q���E���֯/]��jL�]�����.`��Һ�D�ܐF��'�%^%��;z��#�]�.t������iQD�����Ȼ�f��{��Mdp�_�Y��>y�W"�KǬ�����qCڠ2e?�R��X�����ҍ�-Z�ʀx0�f/f��@@�zĆm���t��d�*�� �i��G����X�"��
��Ib�d����"CC��ܐ�N��7��s�2�+���U�������F��c�j��
����H�7Ȧ���+@��h.�Q-�.���9�AP^���bJבN{F���u��Z���J���{�� ��HI��W���l��1��2���F2b�t���|h�bQ��^v�4$�tx�>y�xl���w�ã���v�-��^)�)���f{#�ιL�7����f@� �����a��X�u&d.`�y�����Yٺp�b�cwN1�}RA�����1��$�A�בQT�>fY�y_;�/:�W{(q�/:�T-��+̎�V����-����'=���u�E�������lG���$��X,h��.�&�.��\x1���_`s��� ����`ylZ}�n��g���B�z/�aj��9_m�I��������^�3������P��+S�c��Q�p>�Z��p�ab	/��:	���G_l$�v|P��(�B� �������X�-ºTY�a��o!��)
� �������$�\6$��[ý�#Ep��i%���6(f�ǽ�R:����/~���x��^<�~q푃m�_X��O����M��+��ϝ��׺8�*�dZ�
�"����4$�{T���D�?���BV�l��KK�`�ڝ	��!���R��o$0ۿ&��6������ȡ�^h�$g�_�BOPF��Q0O���AjT���G}���善.<��������EFˎ#��R���?j��������Ydd���������D����R�'�2�:�F/r�u���-4M����H�D]��^naU�ԍ��H<�s��R9"eV4��Un�k��1)B`�*����_Y�@�(��}�����ج>͡D�԰�����e������������ܛ �����v���qP|l?�ȟ���ܟylZ���^@ẛ�R:��`�EB>4%l��u��̱��Ǉ%�FW2�%�����m�����\�Wl/�q$��X�� {>�d2�8ѩ6@:2#D���=�A���st�@G�P�8q�2\C+X�Sd��HS<��?P�8� I�zv��i�����s2�_3�0?����hg�����r5�.y���(Q����\�,�8�ι�V)%��Kϯ	r��TB�h���A �ڧU4r%�X�[+��uH;s�Og�s�A ٨�s>�Nck���aS��]�<���$Zz�X�h�A*H�\�%� 3���%���9VUD��?q�kM�[IĞ������ؚ]�c������h��}��X�PY���%6Gj�=j*��ƻ�W�a+�����n�������e��GX�`�>2|*P*�u���@D;�=l&:w��~	J��g�K��o�,;��i����6���Ѵv��sZ+$P��N�= ̲b`'�& �f�詩�dG�`>�*g�p��-�S���}�q+鶴HզV����&ͣ��uq�MT���D��M�'Lz���?�K�Oo&dsa���~�j�N���D�Fe�[_���N�g�הs�ޔ"�_w��˳[ɘ;���˙vn��|u9��]�T��B�	���SwX?ZG��������z�/�%�=��f��2뒉8��4)K)EY��0B��ͳ��3'�R�4���$��n�Q����x�7T�R�N0����gsZ�s�ǌ�-#��^����R��_�E�׎}����
�1����:؃������Yq�k��N[��Cd��ᘀ�ѭnRw��Fd�3���Kx0��tɈ�����ڶ��0�V^���/ Q�4y�����_.�?濧��'�B1V_��e��ƥf�����b��	'�v�O�\���ܹ�|�6QX�o,����14��z�̐^���}K�i�e��p�1���4�f_h�ۯ�K�Yc�r�����]'2/v�?
#���cј$���������3xj�;ƞh?��� ����:��~�s���7�l|l!��p_}�8��{�i[>�S�.�+�qzL���Aٌ��MYP�A�%��o��9P����q`�Y"*�e���}��̀M^'lF�X�AO�1��8���:bI1iw��\bp1���[,�x3�BѿY��-�A }y2��u��+ 	_  �o/Jgrv� LE�����A����F�.{r	�V�.�ytLri(ݟ[��HԞ-ڟ�|���N5_�e[�k�W.�%�7�B���G����������aA<�;��C�U@���	���v�Gv
zv[Ui��`M۷KU����[����1n��`l�̼7��
�|vm��\i�v8Y�|��	��y"�Q|�W��'��5ܑ8
`&�op���}y�C��������`;XD`s�;Dx�/�[���<=h����h�)��v��R ʦޙ�h��ϑ��*���
���HJ�Z7��m!�5�5�f3�����T��8r�l'�䞬�qE��7�zs0���b�Fs�x��߻v"<�~��T�&�~��8�V��F>�14��4Lg���>>�%Q7�� 6�y�>��:ͳ��.�aA>r��B��K�b#r����WJ�-���.d����qZ���/��S�8����;�	H��Kǘ&��* �����FlB��L|�4�����F��v�I 0)L�~Pې^�\����@O���;��Y���*T5LEW���Ln�	�+�()rOAؠ"gaC;�"�����ˆ��3.Θ���X+9�f�E�����{r�g�`�oJu�(j�a������\T
Ҕ\8#�0�	+F�����5�ߴb��&l��Y�+5�\���r߷>�H�"ݖ�+3n=�N�B,'#�p�H����D��\�X��y]�	��U/�-
��T�j�ˏ�3[�!�E
Ѫ�@�"�W��+���MJ����MT9����ſ��f*;��Y(x>صV�f���T�gt)-[����"|��p<Iv\NQ����3���;P1
Z���.� �l8kȎO����h����*��9��*�����ɢf Ɗ�ql�B���*t=Mᚂq��s`�Nv�E�<0�>׫�4�Xc�F��23r2���vK7��
�nOz�}S�U�A
&�8�,����pq��诳;�	�}�RR]�w����Z��{�nz��r�T�(�P@G#�hTYz��)��3�#g	R����憴"����6�|�v�q*�A�4��"u2��OZv1ى
�EZ	Ѷ�}�����p�H�;8z�]���k�৤	�]u�qa�rl������3�b�~�ײ^8�|&sO�p�!�l�P~`��qS"�tg���y�n��B0���Z��p2'�!Gc��ǂ���}�Z>�r,�PXM�X\�:Lӯ�q(����[��46�Rpt���E��"�
������ {T�
�{ N�G
���Lє7�f��7��e�%��4����'����e._�uv^(�����6+��Pcٞ�wB��k<�9�>U(�ja�c���e�uZ	�Q�`�(,�f�C3?�?�Ay1�7�S���n��.\��_ckR�ME��w��z�}�g��x9�a��w�۠�L:��0U
�[���zھ,	b\���n҇�9��B
vU������ֹ'Rz<_���3���
o [D�X�gV�\:o���hX��m3+���n�j�� Rn֯ESqltN���p��)��H��݊��R5���1mT@���Y�>Dc���l�>�Q�`�����/���{��i�°P�H���gE[;ü�Pw����;x@z
���
��;���������d���w��'����P"�6vr���dp;�����3<��&����� /Ixڃ�@|�R��[>�V(��X���:La�m}_��J���gTԯ?KA�y@�M�s+�B�X��.^�[�#���M������]��LP�[�D��6�L5t�+K�^����RB� sy	�>sH��̦�%�f����+�;��`B��<���@l~�ا�l���B�30�5:Ģf�}�=���Y������`�y�8�0x����k�S��'$�	����ٯwYՖ��()y��T��XT��Z��Q���/	���㗴b���Z|��yNPw1;�^��a�0c{va�b�Za7�dޚ��0�����(G����f��}^�{�U��P�L;/��9������SpH��8��
�^�Rsq��a�M7�$��t��
1���p��8��u���@:/q�E�7+���Y۟M�U��I��拪�Ѿ��'�x�'iо�旣��5����7c� ˮ42\Ð��3S{��^��Fg�j®��ڱ���ߦޞf�f�\
�7H9�A+ZH���S�S~��)�Am��ڔg�s��m�љP>tP���!iմ^uVAzØ��jN3���4��~l˒#};�$����	)����W)$����|"�0�ťɪ��h0��y|W�0|���0��k���z�t�/�g�*�x1ӫ䐷2O���ywX*�v^�p�d�-�?��tU0�5Ka��l�Gxd&S^�����l��*�hӪ��3�)8	�2��yٵ�4��2'���ػ'6 aހ��%]E�e�:�l���*��U��]_nÿe�����S{��얇��?��H_<���#���eUg��^��F�Qqw�t4��� %��+|zn@%�?��6Ӭ����, ��t{Rܭ�+���{�x9� .�����Y0	t���0�H��ĥ��[��s��G	5u9�(D���m�9��E���������u���Fx�����Q���8%��߂�k��K�>ս]K�]n��̆���%�� K��ټ�6S��q(���(Pa����`�CͲ���Y�i���[VJf�
#+��Į̢��J�e�w��Ri��4�.��l��d&�C�:&;��ZES���ZxP�ʢ/�w��((/�u���z�\] я=�K����� �������k��K蕭�`T+�(�����w�b�	�#��|F�O��;���WN�s��H K��(|��vgJ_a&(�M�{~�.}rZ��W��K@�*��>��B��w����v���:�w��<�&�觭��S�a�M�!�tP]Q\��e���sZp���j�.�:��sr�$����^�Տ�>e	�Es a��ZPSn
�3��e��n�J���P�1�Rٰ���5��/��s�@�?�.ᵄ��q����CTD�~��g�aO��>�����)b�`k����Ɛ�U�Np{���p���`�5t��,}��F�!�i�P%�(ՉP�$��o� �Ph{D�Śצ�̚�2�Ԋ1�ɋr��eթ9~��1�O��/� ��@�
��e�Yė�3�U�nN�:.�;���}=�[����b., ΰ�)�:���߀E��B��Ep};Zy���$�P�hru���H�;Np�~��|2:�:):��yk�0�e�4�cr�"n�`�
�Bz����U�$�s�? M
8�hY�և wğ�ה��O;��[�Z�AAV7{{
5D������ �Ty|w�R��4g�,Ű�Y��a:��u}p�Qp�]���!q�,�����s���-4���E�dca�6g��%k��I*�7�P~��u��l]B�?�J�~)�tC9	����j���m�QH�h,��ׂ	��j�?��Y�`��wį�4'a��Q�
j��n�B�#�쩶��SÊ#�����=��u�=e�8o	�y��A;*2�⺀��|
&����0[�;���	�Uf�� T�gaOQ��]����D/�*{qJ���%�l��E<�@�G�z$�D�;����k:=��+�#��C��\�d�76�%I�Z�5s�/�M���k��Q1�R	5˥G*��H=Y^,^�s��W��0PnF�^j���;e?��"��_��enE晥O�5�4��4G�T�^��� ��Vn��J|��U���̟/nG��q������gK�h���+�1�_������r3�9�m������v��A6����Sx��d�C��5*�~�Ϳ�3��f�>�]~M914&�C�������	o�od���F�y��a��zɖ<\�(�_�����	����b	q�fPv�r��*ArEVܿwI�B���@��96�i�z:�cJ�!\�O.��%�N�a f�;��%Q0� �X��*�Q���ȕG�xf8���g��a�Gwz�钼OV�B���-�_�i��nǸ�/�$�v;0f47��j���Z���(SS>�Xx0\������ZD"����ȡm�XQ
�V]a�2�g�7_4m5�� Ia�U���^�I[榩����?�%���	*�*m�g�jA�S�=Z�Dχ���"N.!�E��	U�Z�?gH��u(������`7L�`��b��uT��2��u(�!e�T:��6�c��~a�d]�c��Zè -b�kC	v�Pz�rWPk��[��?�aj1	[���@<���FX*$a�r�Kt�M���(+4gU�-���c�dU����T ��7+���K�o��v���"��>%���<�|���$�kj��k�;(ɳ�۰-?2��`����	}�<�����̼|w*���BoO�ŏ�i�jG�r��~3^�k-�nW52ES/R����ڭ�E���D�'�����|�PVK"�ބ�s���Ʃmq	��\�FFW����$�ځ����^0H�샰�py�n݊�C�r*B���lʚy���m��*�4*�0���S��ˊ����*�&�[78}����`���FjN�Y�%K�����0�ߍ�=�������݅�A�� Q������	Ε�7��rœ�wR�j�K�����7_s�����������Q��A�2��9�r	lq�*�.Lh�{	8Z>�?
]�C����	*?�B�i���kc������bI�y'Ș�]���̄������L 6�S����;�_m���2gnt��F7�i��L��a�歮���/wK��;U澓����1�g �g$��ǯGT�W����jv�V-3�'�:��� o���pր�ul����@���ٴ�!��{3�Q��K5���72GC8~��Bw$GN4�t����GzLG#fvw̋���m(��_���=_ʈ��m�9��Q���b�GG�����bqn
�����R��9�ѳy�ţ�����_u;UJ�l�?���(W�E0��Bg��v�.$������{G6�� �SA5����ZC��kSm8~%+_F�Bio�yn�H��=��Yǔ^�*$�eF����Or ;pL�qG�!{� �{��}�A��i۟Ž�y�A?@E��X<C�����Uɒ[�
I�u^ԅ�we
T74�!� Jw�#�e�n=�f� �d1�p�cݕ����t/�]{8��)�0\��	S_�֑$wH�T�$C�Y��m���w||��F*���a?⥤��JC��:n�º�gNq؂�	��~�`;����3㑆#�n�Np)M��(t]��1Z<���܊�lH��ntjRx�yCh�6�2���Mr��Θ�@i�-8|�Ƚ�6P�̐�|��TxBW�O��o����F6&�<~�F��ũ5�|�@�,�[����MN�Q%d����W�>�\�m�x���ǃ��[��\�Z͍75j�I�1ŪV@BGP�J��_�\��������gqEĒ�V>ib��2��b&@���
[�Sz3�I.Y�v�h��OJ�ո-T���'ŋ:)-y���ô��_jh�����UmV��#��өa�x���A�p3jk�!-w\�ڭ��ߦ>�&E�BC�x:��}�*�ޫ�g�P/�?wX;�K%)n(K���/����Z٣��Q�� ��5^�O�Yj֗��}�\�+ʦ��)	ќ�W"����e����P����<�nc��烴[�F8��&���t<?n�	�_�8��?����H^��z�j�7�q���6�q�e-�q��m��}��Wp[���D���
������B��H�}���Ĺ����w��[#�{��`�he�B"�(��u�U^�;U�\8)e��*��h��%� �V���]�'�-����ڽ'F3��W�����-ΝRjZR�KV���d"�#�[�G�bp��X���pF�fJA���+��ѨEg�;*��6����Q�9����3EO摥-����^�{�P�~|5=��X�}�Y��l��;�D?Ȭ���C"H��L;9��:�s�gh�Ϥƾ�ƺu��-Q�i���v�ȳ��1�*���F�g?��*�*�bf�z����b�_zԋgȗτ�AR�D���� �)��2�����8D�u�d׀�� ���,c\��2�0+G��+ʠ鞛�CG7h��+�1�j``�X^�#����eu�x�8;o;�}�V�_��gL?[�m�1�I&2�\|A��x�,u.�Ga��_��r�d�/��:�q������3n�C�n�Q��G����E��SeeR�*ƭ=����"L�u�#�{o�i�.��ٰ�`/�O#2C����4���B'^a�vD
�׭!��bOb��+ww�� =?5/�k��R��9��)<��B,˷{p���\m�E�	����:���A�Vw0?_#�B}U���u��h���������z���L���n���K�VSq����h�R��+'hu[�q LMV�-���/kJ�����pZ�dNY-v[w/
oR	�7������V�&N`��x.�\� �PN)�$��m��0����=z�zъp�
�-=�2:1&�D�Π�2��f�Q���b�pC�R���6��g^^� X�@ �9��PQ�e�(���D�y�_E}���Ҭ@p7�~ɞg.��@��B�����p�N'� ��`��w�W�T�b֣�S��D/�h)0`H���::���Tf�s��;f}��[:��T�SdJ�GOk��#��S_��%t�E�RY�l��=P�&���kd[�	Sm=Xn���Ƽ}9�bE���#� j6��e��sX�Q��Gv���>��T�Ʃ�--�h�i�d�m<���Ca鍃J�	3Eуbp��k]Q����<t�
I6b���9��_S��'���24���7wY��KE�2T��c�n�j	�y$O�L��z���=������i�N��n�jv�l�ut��~�z'q�L��Dk��g��*�	W��z�s;S�v���$�E�B&�*������,A�.T��O3���p�z�*���É�g$3l
;*���2�K��}�ɛ$�u�qǺT�mA�E��W��j�e��F����/�u�_���&sB,¤�a�b�}��u)Օ�G�}(tlP�]��B�:�@�vk�h���I�+��� tCH"K!�}��	�5�3��M5s����}s�.2�C�V���N��K�@��y�_~��['{\>���)F\�n�'�|נc�x����!Uɷ�3�d�]K{��kI&�#W4��Z���b�]��F��5���16��c�����=���~2��odL!-c�Jk`T�q �zߒR��=C٫�E�(w���/},|93,1�����8�o�D݊�=�y6��"��ޘ��۵Cd+
W��7�h<���V�8�����.U����[Iʜ{vUDJ�}��%�ȍ����r������0��1o��LT��Sb���F���@Ν<�kWnaj��{Pp�5Z�h�*��g\9���L�c�ɕ�R ���¬1�ۈx�Ȋ�^�	�3���2�����o�x�~`�]7��)���F�Z����׼�>5�i]���t-�3(��r��������Zs��t��ǌB˿�UuvZZ�6]��\���w���Q�%��gO'k�}#��̗���z̎5K��1ADO㚾�`iم�\F�q�7��X"r�gx۠��5	z�_Hk(���"@���3��pl��Sk�K�x��%�A
]N*��y�r�'�cF��|������T2�� �UYB�c�_��&l��=�?Y�e(������(�u�����Qf����@K*�w��,'��&s�]=�L/+J�h�If�i��R&O.�e����3���^���O�R}�|:b�7p*��B��c8�z�\�.@�*5��)>{����|@����x]@b��V=����qx�AZ��%���,��&�����`m�:���XPH�����5Y!��@@��/Ob�v�j���6��}��F�O- �hP6��2���페A�%���B��P���&���Lh�k9��EW!��4����?W�P��?E{~���q�C}qL���R��d���-[SC��u��#�z�Ag�i��}V�V��m�d�5T��Td��"�sbϾ~?�� ���2�WF>�J; L�h3����������;�+pe�?��uA��WF;�b���+�?9J1�����Fj�NY�[�f��tc���1U�'�;_bA�J�˫�b^-��k(aV���C"�q������VĹ�ߎC �yЎ�j�|����Q���;�9l�?�B�)�<ץbX����rd�[��7Q�h	�H���d�Sl�jc�S�A, e�g\(1��n��lspu.p&Iex:qr+���-��r���y������{u�ǉ0=�Ȏ�`|zOF4Y�˓�y�&/KP�3&4����:) �����#�f+1�W`S����iq�H���u�1g�ཻ�a���ѽb~��-���"zMo�	��0[�hs�G�&�l�i8j�d�ⵯ��@�D�#��<�W9��"����,�Cմŝ&-heezZ%O2��Ǝ��ݕ]�	�]�5U饁ph�]�[��#�y��j��|W�3�~����@,M(�(��k4UHMe�y�d �2�{f�`�p1M�fw���Z�mӐu��2&v�a�ȡw��8Q�t���
�/���'A��I��/�嗬.�*�Q����f���i�;���s�������l	��HR+/��<`��V�8�P�\�;��z�3��8%�J�6ֻ%��5uR`|��Fje�oV%�|�1����IB@�])
��I�g]t�����h[/m�*������5��PdȰni�%6�`!�Ug��zt�@iW��mP�Iu�yܯ�%/��&k�lb&�9���MGq����`.�>�TJ�����[�����"L����h �6�A�y��X�V]W�E"���~Z�^Y|��;oń�b8�0�gZ����K����_���#$�_LT]2�U���l�G��*pǎH�y!L#�:���6q.���!��-]�A��x�Gٽ!��{�SDq`jf�HF8��8&;��d�HƘ�0K_ ��VOa���4I���;���M�L������XI���W�e8)�<�\٠��$Ujɜ���.X���ә;�g�(3�<4�~`o��\�Г~��Ӝ�WƓ9�׈�z_#��q��7�l8��*_F�Y�p� �l��'��*��
<�"IiZ���R�	UX��/}���H�x�B��J�B���	G���4H2�����C��n�;TP��\.%Of�}�IE�R�h���rK�*�r`�L���0�-���#��������͍w7c�&�H�y�JO��W�o�3%Ufew(�x7�U|z��H���aEdR�����l�_?��M{G�L@�8���rsE7hTnE�+i�OV7^�i���M=w|�	�&6۫���Ƨ�աs�:����0�$X����vA�"��6?';>���<��g3�=�a�U���Ӆ4k� ��j��}F^ZA��eE[��F���D ��` B�h�� <�C6F��ȑ�J��
��A��E�܀�&7%X;zW����+���M�}�U$ǩt�������C�W�ў��1�8'����w<��FZd��d A��na|`]�^w���@�V�JS�tC
G|ٸ��kQ���o���K73c��@A�e������-������V�Eq��b��*���N�NzV,���͎��@h���c�jeV�ff�D@��4�Yi8�/�,le��"wH6�2��a�"q��X�Sa�űG��z��&�jf���b}��=Uo��,��}$�of���w�;%a�5(ֺ9���6��Fr4X:�w���T��3�������'��x	�/_�1����$ٛ�ն=��8�v1�q裧����Ó]�i�C!�GH�ؕ�S������b��Lh�a��@EU?6�i/!����B��D��tI�
��Ik'Ӕ_��1H���eH��i3�Tx �ꭑ�1,�^��>`g�O�9�%�a�`�^2�CYF�}�,����������8����y��u��gfcv�W�7��I��h�zXo��o�D��sfB"�b�<���#�S��t_��] ������F4�l/��h��X'C���	��%n�����'���XhB��(��ZFFǋ0K���'��)7g��щ8�S��c��j�7a����B<��������Ȕ�=��x^ֶ��rzt7'��nݎxt�	`Y�"������'��n������c�A���eK��#����S�.��ؿ�@?��4�ثV^�-8u�0Z]�zH�m،�v㙖E���6�JN+�K���~�����+��-.���m�6�6��̀�"���b�iHÙv�A+���`T������D���
�՘i���u�?�0UN�+�B`�DQȇt��{M���/�K���h���P�6c�͔���Ϩ�*��w/�,Z��G��'�^d"*�f��y)��L�ׇ�կ��-��mİ
�%�.�49ztFF��Z�0��� ��'��1�=B1n���D薂����0�.�A��L�  2�g���<��ȲAK��.}tΑǉ����*6��w8���7m HG�FO��6����0%>`���\&�n��W	�Vƀ�p�QRl�3��Qr�wJ�E�C�	���{���@�D�}r���?�+�$6�U�j�njh>ț��0�M�`�*~������<L��>P�m�]L�/���M���݃�r�\Z�U�����=r|N����X Lm� � j�̩t���3����9��Ξ�~�U��@t��>�q�׷��������G~�&�顗E��	d����
����'l�����%�削�w��k�⺸�4À�<�f��諾��C�'��췖�!�u���� c�M�N�v�ܿ戬���:x ��÷�a&V�7<H��R�=�c{�N�4w���v�P%Kv��e>��Y?�)�!�t��L�u~����s-�����[0xlM	��u�KC-�۹aإ��\�� ?g2<睤�\�����.�bt�d�n4�~�4y=�	�l���)p�3cjQ�>�����ߚ�����q�X�i6���wKҥ�b�@ȭ��'�80\�夲J��p g�z$��Wt����~��4�e�}HDޗ2��uq�B�/��3a&Gy��"4��}��/a���eg���w�[���=�fb\����-�;�.E��
�#�y��Ro���C�N`4�l��-|u[49M�ӑ����1,�&�F�ݏ(d�auW��������ۇ/��)��u�8;�����֟>���2Z�:�,G�a":�}�l�ɟ�9U
��Z^�S�T#~�Y{��^F�ʃ��WH
9&��ױ=?�x���s�<O��U�S�!�N�t�}M���7�&6e�8**0J��tC��y����%�*���$΍�Ep҆�35��a�9]��
�6_E_�
m����%��pԿƶ\^���~UYC���d+��O�k�I��#�L��oE��ma0�d���S�̄'�KP���!
�.]G��2),��Ƒ���Pv�*�_~����M�m~�~�û�,��6�D�be�SI��u_k;�Z<��IoWQ!�J%�o��x]�fH���
;F0����5��4p���i�����:���j��1a�T$Gy9I�*a�CM��a���r�M��5P������"���4��^��IhC~Fp�hF[ܣ(����Ze'�Hp�z�%ag�ǫ9����L�2��_��A.#Mrc�I_�v�����Q6ۻh9f1Q~���fI��Q�DN^@N�7K�VQ�w*�zL*C�4�g$XbB��AZ����jɥ�İb|��E�`��P_P�Jp����>׊j�#mL�/�x�,B���G1z�n~j�l��}�R��+�{�X&�{A�ݹ�,�ٵ4ѓbrB*�Ke�ټ�h)@#���Q��H�oW9m��R�0G��Nh��ٟB��2k	�%�M�`�Y��{����G��Ꝿ��	��X`㺢��"��37Ǝ���k}}EX۶�"����]n}9Ձ7ٹ ��ʮE$yE�R8���L=�޳��J�dK�5�t��Z�vR\�7te��})�]�SY�?� Y��^H��3���������}�<LԽv/C/4!�����\n�����wq�?}�)|mM@���h�ѧ��˄�g��2t��7���O�t�o2��D���Vh�q�v��F#S���Td[<�����%P���2��f(
��zh��Âߏ��?�oQ�F؎����vZ����[��^ �7��1u<�DF�X=�T2�ұ�Ъ��Tn=���{���s'��y�Ý'�4#�&��A���o�3^� Tu$��cV�ȹ|�[(�V �?�9���ȯ���a���/-�n��.pE�6�4�7�>���V��$�Q˵��Y�C`�������w��*R[�#!�,����(Y=�q~���k��}���Mf���'�AS42غ�c��84�yOߨ��]�^�QU��d�ZP�g�Z܊;��6�*=��E�.�W�-���@�mCv, �D�:_�����!�$@�Ѓ�wo����8|��(�|��3-��®-��1�x�Yr�!yѪ�Y�XЎ�O$�����_�����9�`v"����5�P%t�ᖒ�����&��#��/m�7�P�:�q������r�O+aR��vb_CW�V�����a��E<j�VY=6id��TƄ��~F�χ4b���AΟ����K�^/Қ�ezz����S]�6䀵 �6�Q�/�hU�ő���mg�z|����~�8�6��n��B��VG�#����C����v�I.�z;�0�K�T��ڶ�3�8��OP$��h�*��wF� ��)=�P�׻ ��J��5V}?�����X�bEP�H�Y�Ɏ���d�9*�0�䴊�yJ;b��[��_� 4�iY�*Z��oK)�(�@����L0�DgN)H���2�<s�a<6<�$�����h�w�
F�d��G׭$j�_;J��~@�s%(^�x�o�����*���
�����1��8x��o"{�n������]ZcмIipc��W��|UY}��q���$�^{�_��D^.���?-#%'�]1B���qH1���mhIK������?^�q�t����u���%�~�V��[��?ݙ'm7�M��l��]��̏��8i��d�X��^��������+�\���y����h��dǜ����-�Okq�~������o
��|d�U��c׋�T.�'��a�?H�U�<�
�+\�Ą��9(4F�����q)��,bŻر8Wv����*{�
[�f���Q�]�{�m-�Y���/@����p���䣖)�[Wy8��N�W����}n�4[;u&"3�[�b���r���`8(�ݑR������b
�h�W SO&�s#g(�	��LG�8u�=d�@{�O�U2N�V��i8���+�*4��B"j�����%���I���R���%��t�Y�1s	_w),�7�ɬ)����0�A�� �#�9^g�r�P�2�����F2���m� �?�;X��c ��툚� imTY;-�C):7�!��7�������{X¼~&�P��Q����Ǘ�H�5K}!*�K�5��~}����fc�>��lԲ��y�U�	<�	��I��������I&kOL��v��&d��`"h�
�ϹBȷ�i/���mNY�t��꼨�[����V�.�fb��ЂO��<_��8��$^�.]k������B�H�����U�)�JZծ����[N��g�Y(�A<���*	�8��0�j<������U��΍F����f�/dNo B&`v.�
#��#t������.7,M��oQ}��DD��6�\���a��ho���k�K=��C̚�υѲ&�̳�� ��0P'Oh�����U����K<�+Vҡ3	���<��[ ���ʃ��@�f�Y��e�BUy���i�#����#�?B���i��N֎��bw<���M���w�m�U�~�>���g����� ���'�f	3��V(�{��[��1�.���\�^��:����4{��y��p��s�Xɽ�5���i�j����i�����k�N^}oV
��ՈF��� �(��h�7IH݉���	j{� 5��#zӄ�����`,��Gߺ��+��B�Y1v$؏���4�� ���Z�����mys�į�4�Y,��KF��+9����POHy�"��棲m��͍����U������kg{������MT�tS��N�^�Z+�s���ɭ������t����&�o.��'�Q���\p:�}FԢ���S�CM�ޘm1��q6�g2��½ȫ<S基8�D��#	$ie��n��D���5�WE�U/����B{��U��e����˴IO��`(�*`�����_��.�s��F�lP��WV1M�~��<��&lF.�+@s����r/��<o�`��,wL��"�����M��V������=4��.�~5�uKGLP.���/�n�� 7i&�O*�C���.���3��v`���J�zy:�4��?Kz%�����Դamu~Ew~��Z�� @�M��}s�w�%��q�[�]�N{���%�M��ph���W�X��T`�:���s�h�TI��(��%
-������{m J��|��wSx<
�v������_�"���m~Ň7�g���Y��DzO�l���~���-낁�7� ܣX�]X�)V[�-�������U�(eV�K�Xm�.��?�Z�[u��X��/C�cB����c�H���q�
gB��U�>#�lf�J�i|P1|4J`�J�Yh�9���҉w���%?���ot|�@�B\e��({Л� �V�֗>|�cRs����g�1�O@�-10GY7��^��� �뷺�!ܜ��	B���X'���i(BD���X�2�GX�
]��E {��#�����q���b�Y�2{�8��Z�l���6E"�A5�;Z���:x#(w5	3�D��j�͵Z�k��0�WI� ��7�G�Ƀr���Q��i��5�R������"&��
1�������̟�}�Yi�b�Xt]F����<�èud�Z���/!��&m����~28�������w�D-�K�/C�Hň��}�ER{e�Dǜ�!���
R�f��̟֔A�yk�9�z}@��:'�-��<��@H�`��J�=�3Y�<���eE9J1��vr�Wz����E+z�{�igŁ(�8�s<~�ν4��Yz�Gْ���0-�!u�q��c�kh�*��`�pt+��ԤX��D���0��Ѧ���������U�S�WJ�h�q�1��ْF���'���n}��������V�z�-
��C����[d�y�?̤/gF��w`���v˪�zXE�O[s���7��q����@U��r���ǲDL���(f��.���E��x�=���~J����̠d�n0�i�J���0 8��=n`EH��;�>�4���SHո�(�#I�и�/�ϲ0Alaq�R����b�7�*PP��<Z��e� _�R��Ɯ�kI�#��o�gb{��Ӌ[�^������q=��d���r�{Q�ԟ�I�~f�r�S;�_�3�8�|����G��爹��v��*/���Nj~���1��!���#l. ��ou�z�Iȁ͖�<=�9�v�܀�Λ��|����)�ګ ��+������G�*Z��	�e\��Z_��C�� �$w,���h�S�H ��W�.��$���r�-�y6��Q�����n��\����g�U-�e�vw��A�8��P�����3c�+6V]9��}�A|���Ŕ��m!��n���o0��r�0Ѡ�����;*�.���v*`U=�V��<�G�I���P��u&��� ġ�t��|a�NRS�~���P���v�o�L E�9�;�@K���<�]��+o#|KA+�Z����|2`Ȃ&�C���$�x2o� lg�3n�p��1�g��/A��0lbZF���l�t�~�em/.���!�o#����EOz+��@�2t���_��^�p��Ub��sx��cƎ�I�!�<)-�g�D(]�(f;��`7m�ر棰Н��Sꛖ9�Y+M��#/85E,vdP�e���ֈ�]㝘�{����O�^Q�*ۭ.5�g�j1g�Kt�?F���J	�u[萭=@�
���<�F�Q�u	�;����,���N��W�PY/�MBx����f,�V�mk�+��fe�����L Qٶ�7p
O��&��@_���o��i�����ݥ���h>rx��5L�@!&��..���Hڅ8�J�B;���U�w��;���w�9�{�fB�G�U�N�(kFc���'nk#ܺL_���yj��GP�~e`l]$wнBu%�S޲�nR�F���&�bƤ>���St�����������"I+=�b�&�1��G4���#�@���n���6�1B�;�C�ļ�+�5��q���w��8ߡ2S{f@2�Z)fKgt�I������+B@0�^�m![�v}彮dP=�y�J�b�!lO�3��O9�t����̎�i� �+h�a�s¿[@1:"}Z�����̺�h��ƞ0�`b9q}��+�&Հ�U���R�=k�'h���R�B�ʸx#h��J<J��<�
6�N��)ůSd}uE/������Q�a���w�����GG��9�����m�nr�#wŨ��J�*�+�&⹈��:�u%�S� mY|�=z���������|�Ȍ�Ò�@��$K^)�<B�U� C�K B�$F�Y!��p����P� �կ/9�H�<B!�w�2�?O��*1��g:��m���=O
?+n�mEs��NK��(:g$\/֊�x4R=z±��jM���($<��2j~�W.��j�Wk�e�á��R*��E���߁	
I��
��9^T��P��n�e�������?�~5UN)��M~m�?��#�	o@m�˕�h6�����hY�X�d�K�<����i��_���iT�����c�/�����g���Gچ�p��
4;?-���Z6�Y!�	�F��s�)$3�}T�����LNR�b��5�ܐ�l�Y41I�`nס3r������WY׀�ҕ�Q�z<�4�:H�s��8�TB��&��X	\{o�1�� �8�A&��>�6��c��Y�V3١�/;�^2� F�wyZ�#���"�ǔ��eS�Y� �����"|��o��8��p���4����.Z���&O�wCM~��hO�~4�m�d;���ԋ��_�v�u4Kr�i ��ˍ}�`�F�U�dml[���L ��@+P�K�)�қêG$DB�s�}9=�PPl�Eć-�0I�3�������.7eIԁ�/�Qe�&�����]_G����b��C�⪎䋋�"�h�?Ǌ����S��/UlX�x����G��zq���锎NO��#���������m뤇�)*�V'*!��0.Z�8X;P.zw�{���f|ז�~	W3��#1�-�_p�*�.xSO�E�F�Փ�l���zk�-z����9�I9k� ���M�.8G�Γ�_�=R�4��~^��:�=�n]�t=\�[�/M���Cs�pÌ�ᭋ�L8�,,�>�n��s�jzU*r
�|���?��`�А��j7�"G��T�v`���C���x]k��E�
��.�
����L�WI��K�c4����#J4+��"g��Ao����h���4����h0}�e ���JT��J2��`Ywsx_��Г
]�#��\�s�q@z�+	���}�[MᬿV[�"R���n���}�9��"���\V��y�7����=?2h�?/��S�*}�䘻�b���Ob������!���8x
��wl�x#��KbkW2�@�T".Y�%KfT9��e�:�7�K�m�ߒj>rE�1���J�B�a�n�2zV�;�lE��ԭӎ?:�wg�xz�P�+6�N���ʞ�05�'4a��z��b6�����E3�l�T�T�3���F��S��Ȫ���o���F"i�^��h��Q�f"���X����R�]�Y�lG�[�"��XE�J��*�����:��Q	��Uaw�è¯�1���ґ?�` jx�*�g#��3��PI�� s�!�;¾�T��&�$�llSuʴ�ښ��=?��{�$r�ޟ�����&�z&G�n%Ɓ� �Ɓ2)o炤�4ΰ�5�;�EުPr�Mo�i�'�� ��P��|-��$qrv`=�ah�]x"�o�/4�[Rx�����B1�$�ujs����_D�vV�b@	����>�����Ia�5%��-`v�3��ND�-��� ����eçC���<�웥�&r���g4�ެ{��5}�e��B��@���l����f�V?P�6�_�A�����oQ��y-�}�%ᑛ#y�ٵ����6��|�I�uYjaRQ�PqM�N��K���{6�?�/Z��=↴^�@7���F���ؔF��g
3%`	�Aa�vh�!��l��_jC����
6�@�fX�92�u�~�"�m:�ܮwz�s1��Nk�*WnmG���u{�F��L�TՏO	�LR$��8�ɛ*P5�vPLd�xZ���ΰ$r�\���9�G��[F+��Jܻ�I�nx��$�l��a� ���?W���{b� AQn��o�}fԖu���h˰�b���O߆������@��H��B�9N���g�b�o����fr`�Ѧ�ʊA!}0l3�Q\k��l�&Hkޕ�kͿ��8tl;�5!q�B����^W�ƫ���\��T]��7�\JKO�ۍlk%
*̠��A�����{.Q��a�g'@�=x��y��6U�ۯr�v66��3�8iix�Α�����eR�>R�Ò��5w^�_d��wM)�z��~x*��Ra=��M��29Y>MOFQ<l�>�*��)Y+��|r��
`^_?F�?�Ԙ��:��XЉX����	~N��;�vQ���*��Jq.��O�6�8^�_@CH����	���J�+8}jK��4�i���x�����R�о'�|$i��>
������D}����K��*�7�Uz��B�J��uP����c���r.&�U�Oq�'
��W�z)����~aϔ��H
e��j�2Ϊ�J�W���yW����e���;�͈�W����Q�F�sDF��Q�����C��b���ө�MZ���"b�qY-@�2�Gy��A�g9i�,զ$���3����hI(�3	����\�����s^�=0l9��+���d��s
�S�!��?��XE>���$~D侹����3d9���37�7|hm�bܣ�ME��G#��S����p
�������**���E\��/�D� ��V�=�∡r.��)[YQ>�ֲ���P���g���w� J�RC����K�C���g�k�4��3y؅�$�N��%D.d�GO�w����k�J�D��)K�K�Pd���|1��ޥ������{v��#A��	���8��"��d�1A��ׄzU^��R (��Uf�X`̌�\wN�W�B�	��� ��y��r<RQ��a]�>���s��^����5g�~��p��YaكLx�l]������yZ��D��mm�	��F�#�9�c�j��X(̫�t��ʩ��������tD���k��S_� �f�WS�e)�T�~L�D~�:��̼]V�zz�z|���6�2���M��ԯ?�7�п�Ӝ�pz�ձ��	��0*�������h�/�V��'�t�&���C�5#���V��=����H�\���_�,%��b�Z`��Z�����1H�4�Cò��+����»DV�Ƨʖ�RŐM�G�}W9:.{��|[6����4z�T�+u�5��K�Nn䴉p�'�)����ȭ ����}gl��H�V��2��Ǿ��|�� �_�ȴ�Փ ��[ Bع��X�I]��xQzʳd���}���)�2�������%Jd�S�p�__�L��@�`dH(8�=t�:�k��tY�X�6��fzH�J�d>hԿz�D5�Z:��q�l� mN��<#��ׁLk�G�B�3�������� ��ec�"j�=k*�H�f�����$�����]��CIcAv뛳f\>I���lj�R��I��� u��R�~�v�Q�:R�u�D�]�ө%=IM%#��̝P�������sU#q���Ej��"~��\.	�3��78������\.�sO�'�pD�^���5B��y���/�LZ�b���ub��
,�� u�*�~��c�a��*�N�JV����U��s�}�m'�`��)m�\!ڕgҏ�Z!��^KbC�s�fHc�fs��xPF����,����:�O4��	�*7~J�k'�sEO4\ՙih:k.�O�'����$���p�r�M\��v�{����Vt��:��ڈ��� �n�m4(�Aغ����w��g�����y��;b��滚W6;>7��F^��I�CQ�W6�_�i�;u��J���ŧ��Q/�$�֥����|��W�\ʍ����:�.Q���Ȃ��z&ѐ�y�#$�^a��4Q_v��߳�<��g�6c�'���5A����j�'�2�  ��²����73�!��C��Nck����E}���;�c�j�a��T򲂷I��b`���t%���}E˔E�䇷V�F,8�G4���Gy"�z=>���_����������]Ζ9����_�wT�h��28�53*�|�ޟy�qc�"!}l����ǖ4�13������8����. F��[������*�MA��4A����|��3d��7.z7��������yM�A��k�D`4A4.�NK��/�Y2��f��
�K�#0m�v��Q�S��������c0�	�d\����Y��6D]zΎ}��@җW�p��o�@PD��@(HL�)�`T[n?9���.��֨���S?�xl���#)�qo��p	�[]�ݰ�<&��vm��{��?O�r+�f�^�	�{��/�Z<"|SV��,RHQ�{UJqi#HI�R���
��1���H�m��p�H���u�3����S	�nEb�ݯ���(�͌*k���."z�������uR��Ӎ-a-�ϋ���]6�t�9'3�_���g%�[�n��H�"���n��rw�$Ÿ*ȣ>	��xJO��>I��c3ԛ�60�J6�ȃw!�I|�B��Ԗ��R)�=ʥ��K����E<��Nb�8zqZ�]�[b����Tp7:���(R��`g�ԚL�hmf+j�������Fŗf��M=���k����cI��]C{�:Z)-Y�=Hej`�����N_&?/.L#�֌���jq�����~��+&
�6�Ў4��Y�h�4� (s0 ʌ":���G}_����Z����I_�Q�7�mѽ�%�π�aD�6�y��g|���0[���$$fFW�b[�GM,�'��V�Y�v)�W*]��k�b�T�Kޔ?Ć��8/m��� ��Xz���K�L�����J���x�R��:�nD��z^IC�{���u*�t�rx���n�y%�� S<�37�뷱��i��#�HZ���RC�4��Q~!��E�I����;�Ƹ-���Š����#��;��'�6���c��&[1C	cJ{�^ś*�z�Xߜ�8ؤ�>*�iVD��'uĚXjG)գ�|V<E>��X��}��ؗ}�-�9'>[p��^������Vvx��y$��2�:�sy K��֍y`�o�hέ�qxFK��CI���+�Jy�küdY��>��vJ���r�������-����Hu#d�>Z�w�g�b{NК�~BQ3��W��k������=�xJuZ�b#�!���:�]�AF�R���C�9>T��M����}�Q�@�0������م!���r�{��J�NE@����^�u��9m�c��%����isj�cȓz�m��G��E�ZO����/d�{IYX�y��� a��Ib��QZͫ��֠�.���X�W���[�m%x=0%�_K�*�R�aG��o�������i� �+Q�����#^�2�=?�8��t�nGGU%�m����G�0�UDYtu�^��Z�Y'�ڳ3��k����~���=�欓���� 3������c��j�_�2>�JWM ��HV�g׫k��ϳ7e��6>(�MS�8��t��a-|L��{қ6�ݬ��M�U��F�R� �t����?J�ؔ��A�g�� �q�]@d���P�	�Y���1�I��c�h���G��,i1�[���@��{�w���9����5�C�����}��^R����g���/Ӗ}�U-�{H��}��u�g�}=@H�D:���zK,�#�^J2;e/�B��L#�Ak��q��ؒ��ll�&���=Cv�'u�_�߈�<RlT2�|�� n6������S�ȸ�-��H�]\Kٚ-�N>Ĭ� Fh�k|߉0��~,U�T�޽=���䅬 �T,;�g	c3���=H��=hUf���=�aB4OD��!G��r�tȕ��/���ާ�X�����a�����l�^b.#��
���~v9�7���YY��K�:�OH�%���f��Bŋ� �?��v�e����h>OX]��q �d���	�uL-�9�Ϡ�#y*|h�+�WH]��؍��dv�F��B!�DN�+oxx��m��0��t�p��|Nw�iQ���_��}u�2$��
S�!u���Xl1H�ɡ��xa���~<QH$�S�	%�o����T���h+�
X�յ�Z,���8W�ON���4/X�N:��$��"FC���[v�*wD���V%�-�Տ-��&��].�Ev�6+��STN�E9��6�kEB�0����f��H��c��K�	�+����|�q-r���� �jjFg��1켅W؜�s���Z��� �\�3�g�Vҩ�P;gX��Y�<�F�2b�B�a���9��
�S�6�IG�B�5�(I���BLc4?ѹ%$ڏ Ԉ ��9���~͞���o���Q.ol�������|-P������UD��x̡ܪR�z�j�Z�=�Y!��PUQ&0����I��f̱�Yc�h����� R�-�"�+k$6��3�ݱ[�S�/�ĘCe ���ـ����P���]=&S�6;j���=v�Tޘ10�=n^?��P�t'm�b��,��O�E[��D5i��Wa�I�_Hb��%��j��S3<�._cZ.��ߠ���>��o�6MV�.g���l�S�|n�]�M�;9?��#��k/�Z��F�o~��<�Z,0��$z�p"d��E��91�#z��
V%�����_ve���+_�ΰ������_G�	g�}cIH��	�p�E�OlTlq�t�Ȁ�O����xE���j�W�Q������ٿ(�ofm�Z|c���\MΜ�v���	��P�u\��W+�J�F��0e&uj�/$_P�3���rȶ���/E�9�R8��8W�n���h��u254��b�y|j&�L�p߭`�8;��_N=�M�<��7sU��vӇIې�t��,�b����Y����7��1��X�i�\F��>�~�����b�v)���}���a.���3hʬV�.���'��x���k�-��G�����>�(o�sA�̵!�lSʿj���,*7�/;Ef�{����Ƭ�����J����bq���CU�����7l�3\��J�����n
��-��{(d�48+�HWMPc{KO`��K�8����SQ
WC�cW��=_��K��0��q(k�i!�$t��3�!5K�*v$����&C�����e��Kg,?d��Q�4^Z�e�T����L;6Ư{Iu$S&M �6�KڵR딹������m�՗�:!�s�e;5�FbE�|�7�Y�b$WX������
�,�8S����.l���A:��p���Z������3��j.ɧ1_�dڄҍ�g�����OR3��89�������
�
�
�����T���r��(���\��|^��"BB�Z�r;����u�>nt�YK�V��Q��S��X���� �b$�N֐����Cc��e�X�1���?��8�:���2��`?\��^܍��^�}
7�(��^^z�����Z��Ȱ:�ۺ�^f���횒��)<�@I��P~k�8o�����C�p#�B4+���V;k�-����0,��uŃT����Qn�Y�`C�G���Z�~d�bs��p�J��x�pK�U�,`
���l�¨�Ta1�_�*xE�ag��O gq�"���~`Sܓlͻ�6�a��Z�4��օn�6�b}ɼ����3��SFcGQ�Ƅf������z�l�F�a�&o�oV�k-��:�:m)HQ[������=��~����
_;;{7� ��$���6�/�^l��� ƶ��b���UW�n��;�Z&��@�֦�$� �8�E>���V��y�@)f�\$��}GT�
2���}{��O�>Wv��NW���n�x�I��|]�x�>iJ�.e�p��@����_�lfuh��]�i�j�J}Oj{}|�3��ٕ�k�1Ｈ�R����%�:
\�u>���k���Lz\Ii"��U��B��� �W$���^��˙f��9�@��j��W�xyLS~B�{��� �����^u{6��0Glc:�R�#�.�^4����i��/⯃���׬R�H��y�ڇ����/�\�����%2H��⇑i��)�֓���� >�X���x؂3�h����ѭC�e��O��F��N������O��>E+	{�;��Z�&�v������R>�v�޾] u��*�~R����l�+��,"=��5��#g���`HX>VhQ[�5˒�f���Q��p�j���6O��J���d��>jm�)kb�Y���$��:�&:�e�c�M9�z�
���ѥ�備���7fS掜�E
Yҿ�~���Ew]�wIgqZ8 _Z_S�.��*K�7���^pmEM �U��X:5(ҐKgo��c[��x��̂I���-FdYX���A0f,�>Y��h��+Hm2�Aci�N�sHd�W2No�zC�L	ZG8j/`/��yؼ�FGP!#�0�j�ndɳvfA�6o��`+g��t����F����l�`5�fp��Ї��w��/`=�
���	��;�W��A0�]��I\ �s�W�<�&r@-"i��=����0�P��5��� R]�1�\�)Q��l��YL�"v�B�h�,[,.�"��;�h�v8�d3�@�.3�	�L�Jj9i[���8�>lF|F�8��n�$��$%���7>iTx[���q	כ���8�n`��6G�)��k���DS��2�x�bvĊձP}����l/��sQ���N�,@"�.n��r,ȅu���j�Uk����PH���ӎ�)��21�Aw�~��g��ye �����ֱ��m0��%֛FIՎ��Hɍ�<��u)	��^��#�0��$&���Mu���*tY��L� 6g3�y���ԵԲ�÷Zڄ>�_7���.g�Q�E=S���3�o*��W����T$�m�8y�B�-8��\#��G+�~B�j�-nw=}��pv9<�Y�~��3��[J��%�`GL	��Zdx']U`H��"��0($T���a��r�-�OR��{4J�^��v��w^�j�,�O���v��~T������r'��-��"�#�5c�J=/<�|��?���l5F�@�<�݋�4�L�m��!�ʕ.��|��u�J�Z&Q^J��D`1Zu3�/ϗ��ܲO�1�Ǌ(�g��q�Ԍ4{���ete&��޳&��E� в#t0��L��.���a����4X��A��=-
.����ug1��س��?�b���lM��b_Hp=.9�A~���,���6��1�l�C���҃n�.t̴�#�2���(�󯆭��=�]��r������S;��z��%ySw��1�/�5(��g49�M������k*jx��i��VD���d���:�2���Q�$fԾr�Y�/Ĝ������|�&�yk�,=�Gpo4� �%�b�A��U>q��`��Tn����Ym~C���TM�*q�Vk�&���fGS?�2U�Ԝ�R�P\��s'E�y�hi pY�@!��y1/Lռq��	F��D{O�fˌ�оD��K�A!����%*�O��#�B�R�ң�\or(!�!VPnG�E���Mv�"�5���]9�*p)��2�dF��q��q9ox���d�W>�W_k�u�6�M�L���������lAᢈ���yA��lk�,Yks�Ҵ�oC��	Kj[���֫��-Ԍ+t�F�e:�Ԭ�I�
w9���� \M_����Ć-��l��I����#�Y̅�i��v+��h�(aM\q�|n�Vvc����z�-*��m]�s��mi۱��0��Kŧ��瀰�.Hǅ�~��^�L&��|����pq�[9 ���ՇxUc��c�6��/��Z��8f8�Kr�]R���0�6_�.V]4v������A�?�^(	����<������v���·�Xm	2���tɉ��}pw�_�Z �r"ӆŁ#�b�)?JI%����lƅ�
����_EI(K���J>��vz������V]6�&##������^���+
�/�\J����N����b���p��-�����9��)K��[�����d ��rv2����ߡųw��QTRd�����C��n{>�U�n���R�1��33N[��CW5�:A�6����p�W�����A�e��(m�����ה˒w�?�No�ސ���wt�Ȫ�gF��h3��s�#�"'�PL���7���	��u�@T����8z�������X���\�5)y�#ɻZ��{"� �q��Q���ȱ2S���Y|P�ջ�uj��j���Пa4��DhD2��T��۵b�v\ ��_���~r�b�%`)����=�|qjh�'C,�[o}jۙ��n.B����WOe:�U��}���{g,&V5#�*d��>�T�"��tA��2[�/�ԛ����Cg�[��$ʻ��K�2��S�W%���"�F�,
4/!��ۈ����f~��%���A��Y~����eݣ��*y�eUV�Xn|;:��(��2&b٩�F����^I��z��l��3�����`�t���q���xs�`V�'Q�N���Q�Y%�ѾĊC�	��������;����/���q����<2�|:��c�ہ�0������z�7���;��L���(���&ZK#�i ���0��j�Nє���7TK��r�ɋ}j8���]Y�&��!6�o
G��ۺE�zQl��>��(�[�Doޖ�M�^;PD���w���W����HOcG�X�Y�}�;$��U�|��W�ޮ�D�'�,�I.q������0��i)�B	O�n���
d�����<���E��xVT�sim�t��U׬��૱m�5�YR��� ��{PV�7���.�c�J�:�$T���+�G݅��.e��O�������VA�{�×< X3*绡d[�*�U�9.s�J��GiX�T����B�����\��x�e�J��Q��X�ND��Q!����BJ��gZ���f�~	��p�Z��ʺ�����e��?��0^�J�3�{roI�uV����߸/�k�uP�X���Bz،b�(�攽ґog0��&���Q ���c�Ɇ7|��GW�)Iz+�Ur���䪱�_]^�\�:���c2�;��K��_��`�QX������X�5�qf�T�Nsǧ�\b���.[�h��F��њ�KfVׄ��+�h'� [�]Y�ߏk��!7��*h}ٱ~\M��$���&�ɴy��+�_�/M�bׯ��t�K�)����K����2{��n��.�1�f<�W���E�?" 
�^&r�L��O�Z�#��C�%We=x�h�0��3���x�O��Q]�<�����
{�V`�2m�t���O�:��P�ÄOs��i��Y)��趤)^�q|&���f����#1��Zv=��-�Op!e��\
��2��Q�r�>������@��Y�
�[je_6�T�5F+K��]��\x4���L=�bN��MG�z'T��\e?= �:>�m�*r�=��|2"�$�7/hW$�/��1�2hq�n49*44��4���a�0�#�u@�R�!Ʀ�<a�v:X����Q��Y!	rgL�`���<uo8rO+V/ m��Rw(�p�3�ό���cω����АM�4RD0�`��%��Ft�o���Lc�&�ɛ�R ._�3�s>����a�9��0�n]C���C�D���e���M�M�қoS��q}�������e�5��Ve�#m�%+/>����͞~��z���7���H
Tv�W���� ��<EY�:����De+�0�"?�����߭��CH�����<�B����fU��T8��WSq^ksm��S!�֓ㄢ2�`����U@�X��M�]��IVBiuN,Y�B���#z�qJ�ݗ�J��5�n%Ux ��Q�D�{Pi��;���6��-/F7��o���6�[��C����4��;�
�|ڦ�l�o����ͻOe��� 6l;�c����(�(y�`����tp���#��Y���n5�)�Ǽ�q^�0���R:��%�a�F|�oG�S��r��A��ú��ׂΑxq���Z��^�n�Y܊����>?��?��U�Gwd|���B�-��T�2�aNK?��^�t�So����I�{�3!�a������p��x=�zz���хV$F��k�����D��i�o�@���g��.L9!5HƵ��txj�U��Df�����������.{�_K��ǔ�}vn,gw\��8�ɏ�zCy������rT��{.�#��r��>�&.�#"�l�X8�l��J;��U��;b�@(Gj�q����(u��e��	���:O��~�˰J{�fva�$�Dj-L5��rk����S,bs'�Ro�tI�Ѳ;��w�a��횚.Zdn慬����<_~w����^j��Y���/���.�al�M�Q��x\a����$��;�����m�V��}D���)�6���`�6[s�����llr:h^��{%��i��$RY���$U���8٦Bw���?���[$�{2*@���ui��ۉǖ#��Q�ؐ�����-2Qɸ)6�.`(Fm�V�i>��T�.�1��q������#B���8�lX�� ¼j�����3����k #�X�*����� Ak��^��)��ɬ�r����s��e�*E�ŮḢW�wt,�̬]��ò�#:}��e(p^k��>Q���Mj{{��]�qM�[T���G�Մ/S��2�q=��: |$�c?.��#�c�C4���c��G��}�Y,#W�B��q!�����h�>��L���HB�R�&Lݵ�p���fI-��+��ҭOS��_�]q�8��=�g���(l�g��/ ��$/1`lK�[�����gy�b�l.U�S�)��7�|^@�r���S�y@B}����P�p�� �f~�1ӿ��G���?��AK'�^������T��s"qץ�i:ގU�F��m�0�X<��BSb"�	q�����@��	��.�."�G��B 	L�`,�q�ʏ�2��+s�?�\�����2cʝ��0.�=�D�Hr��8�CB��e;,��Z۰�I��\i�b�x�~�柽��y֬���mѶ��`Pm|��wD����=A��e�a�dI�&�j35��λ0wsK�9x��S���m�y�tfq��؇�pI�c�?���4����A ���T�� �Agu�9țSw}�[^JT�G��*�eBM(����Bt��H<�)�	���c{�)�3�hs�����ˋ-~DG���	4=��'(�皤�\X��E Ev�ᦰ�iH���e��ǪZ��N����CN��/�BMt�|_9�ۢ����F��ey,�nA�l�'��psfE+t�`p�"�7�t�����V�0�7�y�aI0���[�kX|̴T�n��<�<��MB��N^=	�L�T��ژ�/{m�{��@�/V�8����۝��wW���<�'���ul(Y���������âWO��e-��2&O?�eD��*�~U]�V�IqS��.@��:���ޗm] �,�5��k���*@j?|/�(�� xyA��@�B�!
�I���ނ+�K�V�8FǪDs����NF���LMD�~P1���E���%����t�x�f�Tf��%\�������C6?6W�Ux�kz��#�w�[Ww��u���w��͇�7َ�4t��T1�����!��1v��"m�-|������ �,4��N ��$їop��ws%�;�V�����614_`�|\E��O�ֿs�=:���T#� Jm�+�r<:�!u���<�e��@gY�ebQ�����RP#'&g;��|�v`���\� �ߓ�ҥ�/@�R�bC@Rw���?y�U����cr���Wv�2}�X'֒����۶Aj|\NJ+��O.��Q�m� �z`��:5fK³ϛ���N$H퀒Qߩ���%�@2 H��bX�:D|�v�r�c׬�#�ٻ�-�;$����K������sWWJz$�Z����'���Q�_[�R�[�G����aD.��
y�G�8�����e����+�J�m���^��;9>�1�j���\�}�2?@�p��7[l�P��{�2,GD�H�?|!�ںd�GAu�������	t�?�"�M<��׫�����ZqV��Pؕ\�Tݣ+JYx?yH�h�����W([l-�v�����-����
��§�=��w��w[Bl�^2͉�cޮ�.ї��PXƣ�k��Q��.�	b������|'1���٬k�%�Z�ݓ]�iHԖ��XAH�l���!�eR�JNb��2���Y�.D^Ƙm*�{�g���+�yc*e:�1�(�!���y.���0�����7��W@�~�y({�(�kV���o�f����� ���_p�H��HA/�}P�Ț.{\ICH���C�|�-�R�g���"L�!h��>z��mʈYǡ�=�z���*ҍ%w$�/��c$ ���R�S��rr��g�\"���e����]�=�[�b)�z��V�T�xݦwN��}δI��Yz7�*d���a2�\,e��ŏw��&t5����R�|�����k�~q����PPa�k���r�Q6s�?���G�Hb�<�Cuoć�b�����k��w���&�Z,[
LwGSf�����Q��zŎOTb�%�������R,��990�#O+%�̬j�K�]�V]
[�9���0mc���y��j�A�\�ʈ��}Y��xvCfպ�,h#MRiI�q�< ��y�ņ@o����%2�Q�V��|����c��=����!�I����BN�5Ֆ��S���ַcz�*��Q����#/'؈���x��/�L0���3��n�8�&ئ�.E�:/��3�z�6j��Q���A8�2�E�X_+����rD�e-1U喉��S�`�����P�"a1�Z��؁��d��<qZI�!ǘ������/�/� ��X_g=�U=j��K�- o��%��b�p��L�ʱ�e�J�����wB��j�]���t�(��K�iŨ���W�'���t*����Ph��C7�h�e�-T=���]i����:�6�隧6�X�5�LFFR���\h��g�Y���d��!��#Lu����E�ޛ��G�:�w��Z��-d����0���|����|�D��qr�F�z4�j]�L��r)љ��ӳ<��5�R�G���O��q�����;�o(C%��(�eÄ_NK5'XF�h�`�JZX~��X	>7Z�xͼ&��,�b��N�i������:Q����m�z}��۬���R�D�����%�tmS"���:
-���0c��&�h��>�0�7O��zl�`~���5i�z���V%e�s���e����cI�����L[�o"��W1�� ��~�[���@��x��Dw�O���3 @�u�r��\Ph`B�&^�	��j��$�a���@��g�Wv�F�@}>�sٿ��<m��'U�K��b��0ʛm��|Zޜ��c�۔�^O� �)������k$�=��o�Y�&' E(�:�bQ:�ݑ��26K�v�����>�Z9�3��j�Q�~���z�l��*"c�~�]��s���n&�9ZR� �+���Z��pL>���!ZZ�C�q�<��q��VtD�+��k|C��iσ�]=E��N^<�[dj��v��	��S/{f��|���Jj�<٤IS<������0���~鸸�l�J��7��i�9BTAX�z�`��!��2)Ҹ�E�4i���Y��#��|.)L���dӽ��D҄�.,�d-k�xHޮ]m+�ɶ��b�klR�f_��w�a�}P�|k
1Hr����h
�&�|D��e}���F������!JI����OA��MM��q !R��l��ѿ$��R�.4Hf��2	qJ�04t뫷��gǟ�2t�j���u#*~�6�.�k�e3���@�r0N�
j�0��^�U&c�!�>y:Ȼ��k�`�=��:������=�$��J��c�mR2{#���[XY�*��c�V��t�����?�L�eB�m��e��_����"(՛������5�RPq�x$�?�ȁ�s?�5�=��y�� 8w28�Y�3*ł��}�SA��A��E����T�?=Up1R�,��d](>���Q�~z��Z���������x�6�����/jv?F4���g�З�(��ؠZ� ��7e2P|Z�I����B�.���a�»o�'�^�N<�MROT��(m2�[����a'R���Y_��rr�jP�
R�$Z�J�T�!;����8<�Ȕ	�+ ���tDMT�	P�)��j�9�_a�v��.�tç�'_sȃ
��݋�`�x���A?4ie;!,W"��R�>T�?&����L��@��1�2���{ӼK���<�T��y�P�~	6ى�ט�Fȅ>3�S�D�%.�i��{��X�lt��A�&x�sK��6�pՔU�T#Qfmێ�yc�fv)i��d�>o���m�Uâ��]�V�.��<C<������W��"l���������a8��N������6�y��͎d�����ߣ��&��r�^D}ժ�����J��̷���=ݢ�J��~N:�vND�3I�*�=�+�_�)Ր�T<�\����_2N{r&����i���Ç:���%��ᵋ	?%�ŀ�%�1� E+ H�UH�ޮ{��i�仒��$�4���A��|	Ӽ�٧�����[�W��Q����VI����Y<@	}�`>������)����&���MX�avi�Z�85����.s_Aу�#���BB�oq�ل�f��M�
�B����8�6[�ף �A���<~��O7�<S@��7\�3��W��A6���:S:��;A�����Rӏ.�h��-taϩ1�2Az7���Y�u�.����Y���is��}�kˏ��z��s�<WPj�A����3R%{��+�UZ�)�BW\�ai�Ib'p��
0kz�Hf�/�������1��B3���/n��f�j���T������$G��r q�eY��C�2�>i��dlM?�2֒:�m6��JWoW��k���"�»F'ᶟLį�����sV��b\$��md�lt����'2��a�OSL��m��U��7�o�fh���`j��f�/Ee�t�n����!������7l���l
���YU0��PB�fu�s�����m�σ}b��T���[�e�/5X���I�nEt��es��^�E1��qx���X�p��̟�|'�v��[M_�@(f]z'�_�)wv?
��*kD��^ӭ]Hg��s�[�ʟ��g	��D����C7 �~�`�on�)L����'|�� I�T3ݷ��F�n��D��w�z�t\4�%��Yd- :�X{�Ye�fٷ�2z��3@�,X�x}q�1� -��A���Ʊ��q��_?��H~��ReS�:��&f�t��-�：��@���8uBU(�*-�� Ǧ�-����~���(m�1��lHN���t�#L�0��fIF���ǌ��c4"1���OP���GF嶲hXz�:�Zݐ�>����$�9��$�����7�X�2�#E�����ō�m�9���0MJ@�
795/eސ�Ĳϝ�$�\�)8�]�M�+~���T�1��jeF����/]U��[�7;%vU$���S��ϴ��S:hO�xJ
��X���;*s�2�}bOAb/c�D-�+�2[�r��k�-��j��`ޞ�3w�0�SD�(����=��
*���{[���2T�2'�Br���e���)F��Z�lnv���E�̠<�綠kZ0�P�:�j���?m?�c��@f��[ߠҠ�����(tjsp �nW�!��F�x��9����������/j�Dmg"����>�����O7!����Y����W�N�6�{��$��D��i��h�`ɰ����?���c���q1Kj�E�B�g�	ҁ]ʶH6�*�\�/����]�0�7ﯳʘ�` ���pA��i\�)��>���w|�;�_WU@]�})���'}F�U=	(��G��rE`��"��~�*��"�k��7����{�F'�QI��D"�V���u�������4�����~�¨���ɐSV�T�9S�#x�%�H�e���M��Տ��2�"�_F��.	WB�_��nm�
|*I4���-��� e,G����-��חLA@m�p��m�K��Xz�^���塳��VT�r���ё�A�@1:�c�l�u�!�(�o��b��G+����D���J�P�<�Y����/��q�$Ⱦ�M`�m���7Q��R�f?҆3��{˘���_*sΛL�8��8��\��J�����6�S���YԪxd 6��c�Z�e�,p�7�3��Ji�ۛd[�z.��2۪,Z"�8��tCڶ���[c}��tOĠ��%0H�kT�g�2��Sk���`��S�D�8��|���������P��8!�c8�j�]�����yi���֟f@.Cq�E�6��#5n
��q{�Mmޅ�i���&�6b�00:�g����~���۳vzb�����w�hz=��c���:���E����i~ϸ���tU�����G�a�5�b]������|4q��o�0$��B�v[���.��Go7��#���[��=[�4s�pc-�&�歂�O�ڑ��ۧ�[����T�����4�ib�O�^����;Z��H�Q�1<	���~�)g��6��R�u>sC�#�m�����r?$)?���at_��$b���|�6��<�(�vaSjt�Ў�#���ߩ{bQ��@3�T+�z[��*�S��x�P��`��$�B%��HU]iWW�
~��~Jʛyt��S��"9�i�%&�#�c��������� ����c�<.�'�T�,/��Q����RٝԱХ��
�\v�L��h��!��J`е�_O��a@��~������N���L�dJ��ԧ+W`�``6�Zm|4sn|�ϭycF#�EI^f ���n��$���36�:pK������T�	x���ӕ�g���r)l%x�cI䐰O�c����c�R���V�&ywR�eg�����a����5��Tj������JK���J�����K�"dRZ��&`�i����ru�>�#��	��®34�L��	e�y�В��Cwל֭��k��1��/�d�}N�5y�m�?����2���<���HMѶ�.f���9�EA�Z��Z4�]�^�v!�k�/+��h�Rx�+��oE�%�S�����/S�f�b�俁-�`cH��]ݳ7�Yh��Qܚ(�.n6V�*Wm8�5T�
{3^��֪" ���t�U<��=�d0mH�O�@���"a����,07����0O��(�{;Mٌ����\3�wK(КVy�����F vl� ��Q�����Q�Ǜ�%�lV޷���j�٨�z���Z��6]0�0��B�:\�����O�;���c����%��M�p�)�z�$&���3Fhfyf���BD �_o1FB]�д�yF���K���VH";ɥ���Ó�7�2�x�'�4���H�!�uP��ɞbX'�Qax�\$0v�|����30}���V[7FJ�$�/0���֊�|q���*k�r�J�2>8fn3-��r�w�����孷Ρת=.�8g#&�h��o|�9�}6\�e����a�w�#P��!1�x��؞m�M�s��B���';���KG"��X�x�p��o��"��)��nu�I��m�X�Y	�5���9�bbq7R��.݄;����WDIC��ׂ]J�>~~� ����q=��W�S��\����f눫�,LZ��Q]�q�K]���=-��!��w;J�Hrr�k���nqg���؃L�_�!W��3�j�K�&:�-�jg3�\T�R��#<Qr:��BAX���U��z�nb�		[9��*2+��p�I�%��O��}<<��J��n���;4�.�v�w�^�@s�9��^�|	���8m��H�!UI��8��K;��a��n��(����-x��8d�y��#�źP�Si7�[�TLբ�J[aJ�%~�c����-���yz��ٛX���8-�x�A�>���P$v��yN0�^_�_��M� Y]^q+����͞m��t�BodJT$+oY�'\��sU�B��ӂ��&�(�'�.����o��- ��D����T�N�0���խL�mۊ	��W�G�=`�}T����yA��̊T<�1u�ǏT�q�0��V!`�\zs�+f�X�L�����.�H��G�����9������<l���XuQ#����S�k-H6O� ���_҉B//���QƤ�UH��{S�	x�ʝ�!W"��V3���O��@���g/�i$E�C�38�l���#�h�bfziu
�r.���h�@��8 �����*:B|>3кP�Yvn'�F�>ܔ8Ьz��8Ĉ\�	�|��Po%5&X�� q�x.^�ӏ:��aդ�|�<D4�խ�4cG��>�]�݌���"B�*�s����×ZV*.�W�˫�O}M^�wX�F�ȼC~0�(��72�#o��x9���Q���<�$�� ����7V���	�z�Uذ���0 ��	hұ��ҿ&�{G�JpXË����!�o�7akf�]��w�=ď�dw�=5}m���VfGpf�^$��P�Kk6`�ds����"N5|_���C��;��Bòmi3h|Am�,C��z�*!1�ڞ%�O��~_7��A�)��@C��0K�\�p# z�ჵɑwe�5�}hғ�o�@=bt` 5f��Zl�����Q��ce��T{3,�Q�No϶;`����=���x� ����/g$���ش8�����e�ã7�����KM�j��#�3�e�[v�Y�Z�|=��DZ��ڨ43}M�M�*L�ػ�`!9�����\gNЉ^�A�h3�b=P�9�9}Z斑=�Czic��I�����+bՔ�p�Yw���t:0h ����)ju��Ș��$�p��������Ϯ�vpI���k��!g�#�oC��3A�?۽C;K&�JR�C)�^�
'��>��dn��G��>��x4���
�[M��a5*2A&:S���<pK�cl��+���.����r��c���N8oچ}���6s��Q����|Y��peڣ�=+k�5u�g�|rF���g3�[�\���Xw��8>�|1�"�@���L���Ep"O�����Db�s��F�\�i���]��t5��q�8o�񘒟7S��r��C8^��m�K�r���|�z55��\V�Ѿ��a��k/��r���l�4H��Q�t�o7�ҪV�L���H�E1�m1�Vǹ�S����nXF�,���t���瀩�
��uК���\6�u����N��gh��T�Yf��K����3<�T��<��r38#	u��������
���$��!���$��f,���@����'��B���	og�j����/ψl��P�����,��Lz]o֓�UME��)�c���v��vd�V�A�C]���'���(�"��*^ y�Y~˯GҀV��ى�U�9��?㬈9E�˖�w@�.��+��J`�N��
�gB�[��b�m���u���m��]_L��1�����H��?^]$��,�~�'�'Q����%-W�$*�Y�ﵨ��N�Z��H���O��O;���e��vt@,�8�*3`�X�+%M��~��8�L-�����LɄ�x���\3d��4�	A�a���c�>Aw������eA�:��9���Q�0Ȁ합�����K��������%jB���m}k.U�[���厗�'#,0�|͟�wO���&���_����S1��ؼKZU﫞~������ZS�XsUU
����#A�m�݈�`�q�L�HZOd⦞`��6W�;lV����]#>�i/=2C�/A��eUa��HQѽ�M_c�?�OAp��"
��(����3�r�i�����I��fCY��d�&��a�հ��g�{�ǩSM9GAq	����r���h���"�7�wa�o'3�b������,��h9^-�B�2������i�Ik0=I��y)����[�����T�m�����S��Y�n��jI��0�8M ��l����C���8ƕ�U\^�x6)�8��!#ǭg�D���Y�wN����=��UÞjbf݄�.T��E��a1�9awwVx�����P�� 8��gP�\&���b�>9�3`��j�O��z��Dg��`�j�oB��<�qӧ!{m\F�1�5%n�P[m{K�z�m��0�{�N!I��m�[F�wf��=5"N�����U�{�D�K�y�c��= Yt�b���]xHe�m˳��U�YWTR�ٛX���+/��-�����qN��+NuO2�`��U���O�jա����+I6��y�.Uf���ԅ0Š�� =Xl*���h=x4���:o���Kִ�'S��V]�-���&]�4�Q����0'/�;���J�o��>N�}m���C�����VѰp�y�����9��W�~`�mb�d-��G�'�%rJ�<�`,~l�u�����8���5�O9�Ď�j��l�o����Fii˚��S��Y��d>��R���a����!X}�=b��-f��U7�x���+�R���k J�P^+��}�I�frZ<����X��s�hK��Nc�m�dC�����6��x�4�G|�Qw��/7�n�Tǚ��w���<)�Np��p���r4-ǥs�\okwXf�;ag��{W,ǵ��\�#l2sґ�O�,�q�+��ȡ�A8�=�zQ���ƙ�1m�'�%~����Iz��77�1$�:DĂ�jm���[�5z`�F�ڛ^��A�d�� D�+fM���*Y�܄^p��Ǻ!_޶�w�(E�@&	:hU��-5�������'�J#��2,xԁ*�d��1�:��glV����ӳP���Z;<�v��� ֗�&zZ���n�V�Qӫ����ٕ�(WJӋ?���tL�Aʐ��#���3��	��$px"� �6�1�le ��]�ȫ��֦9�O�� �N��a;G�9�^ �:��&�'^K�)W��UF�893�Dc�����%ZS=�"4�O�������6�����@�z.���ֲǀ0M�&�����ƲXl�ƴ�o:�Z�4�<:ȿV���S�l����]��o��a�>����uW�*qL93�x�S5�AO�߉�Z������#z��$������N�^w��J*�/�&d8�:�x�����RN��= 6vD�UG���v�7O�-	Lel �X�ì�����LF�&L��V?ڪ3 �a��E� ٴa쮸%�H&c�.I�BM0W?DW� 7�`"(K��S��L�� 6:�7�y�F�+2o��99��0R���y��TY��f�%������aN:}5�<Bh0-���N�b�T��c(��X��{������VQ��h	�ni'���g�G�6����G��?�#��?�M��?t[��� ��C���*�v~3�a_�ȉ{�)g��hF��G�[�W1�~~���
�e�5���M��aۑ[��O�̺�[�����u0:d6�EXR�Uƃ��Z��j���F����ʹ��Ww5���D��ŋ�1\�� ����\�2 �#�dj������ep1��95ے����!')qe]�����Kv�e_�E������FsCA��p�m���Sy�N}�&�	�⤾���o�|��z:�
o
���I`Ū��\L[�(�$#��ۊ/�c����e�PI����Va�+�v���M�,L����[��#�����E��`���D�A�	%T_�ݼ���
�����L��̕�δl�mhw����?T!�q4�	TA�o�R��g��a��8�֟͝�8��	"�/�AWx#� ��p"V7�ЂҾ���6�2Vp!Rǣ{3����)�d� �֐��jA�'�h^b�\Dj 6��&�@!���������E�k�.{��0����cIY� �nXAtq,l?��r��?"�(���s��c _�wl�dK�(k,�{nQ�F_���+�S�Z����8c��5��K�m���L��#���nÔhw�IT����Yߢ�d�N��?�1�iv�~riFk��r ިh6QP<����C��e����"���!`Ɔ7̿pC(6�؃N�u4�����Ӡхt>J6�#o"��)cCn=�%{Ի����:��G�8p���f_0iY�o�*$��|�=�F�M�^�D���C�5g�V�ŧJ>]����R
2#����=�����r�a矨/������gB�`�X��M҉8_��o �4g�u^����%��m~��P�9�ʡ�S#���LR�GU?���'ia�/g�D-���r!]�A�b6j�{�3����rzY{o8�kŬc������+n��������9���hl������w�k�
Dfa����w�m��[�T��]������ %�5g=��@����L���zM�86Dou����9�XGŻĭ\/�p�W�}"����z� �b�`��6��J�=Q3l.�zq���+�t*���{�l���k���҃�ct���j����a~�C���t�D-v�#�N#/�^��
%z�O�wB1G&w����R��qim�#�ǽ�wX1�K����:TZ�<c���|�6X��QJ��#.s�:��Q�7Ш��B�?eY�A=Uؘ�C�n�C�D��O�����$��eb@۲@yhj����r�bp���d,^�����|V,%K��,'����b}!3Q�T\���]��@#!���{�AU�������h�{��u
i;�W�3��à�0�n�i�qƆ�F.�⑋/��G�B����ZF=a�f��b��^,F�i��P뼜4��KS����Z*�'W�O%�2t��:��t6�fx<gg��cm�U���aT ��	�s��K�uw���s�Z�mKPc^HSy#f����4P�����}���2�$	"71�:�j�U�)$�!� �
��<��J�_Z�7�O�Kp?9+.��틠}�<m�u�9��ܕ0������d�pS����Ej�ͅ�e"`���9��L����H�� ,���H���׳?�|O�g
�a�N��EL�z˿��i�l�tGGK�c+�Ү}��k��k���ۯZ����x|�__��z�AW"�*�<�\d02�l�mP(�!�ojCX�a����j�E������(Ͼ��ʠz.�\���?ӯ>���ݽ��9�B9���Z�#.����io��=@�=e�D�P��EJ��g�C8&0�U"j�����B�&xK��{J�AL�3n-*�E�`]� ��=#l[��:�.�3�i�:�V��G�I�hBi�˭\���˭��UB��.=�7>�䱝�`N*��vpqk�ac!�	���,�8�l�;�zQ�E�\wЏLϣ���N�K=�x��t#�u����v���B�L8ǥ��F�db	о�C��v \=R���X�0Z�:�Ԇ�:��{}\tAj�Y�a��͚m@��s:��s�<=�1�Bb��r���a�<��f�~���������T������gpt�E�q��j �*�.�)b!���6���/VEo�����Ed~��`y�`67ic�hV�:`��֩� ���I�[�J�\���/m�c~�:�i%8^9R�
7�o^_Pd���8S��I��Y���g�%�W��@"!��e�E��1c�w���d��=�����&T������(��:�&og��a�%�6��9�)Y2I���O^�4�]����fȐ�u"� ��"�.!�Udz'�H͔��������mi1I]l�2B���S�~u1,�O����& ��1������ �'�^I�7+�<@����ߥڨ�_I�=}��obI����?A�v�<��-L]+sL����I�H��eAⅳ���$�c��b�ĳ)	8ʞʳ�{��"|�yz�C�	gH�zm)�������p@Q�ގO�J�R`@l`�r|Ō�n� K������ȢC�1���W��JU�������]���;[��d�K�ɫ��k~UZ3�1�.7�%��A?����ZdX(9e`�\����'�]o��y�&��xŤ�N�GoW0�7B�m+����bhO�+�u4���TDP�[�l�v~9<N�q,���~��tG�߬�v�x'�����4�� �ě������8��q|�qBߚ���?&D5|�+C6��y:P��5E�>�m�}��?4�]���Ya�^�#�P���J�ϥ������&���sc�6�m��OК�,�����l�|j��NO��Nt�����ԡ������5����)������!���]�0v�Jn7U��:��y����`���|z���V��?�G�l��_�"a�y,1Ƿb�A�����{�vD"3ŉ��X#�����3]`_��(&�h���w�dƚ*� McP.w��mk����Hf�wI�Zo�$�%$��S�k����:������@�|�T)9�!I�8���D���m��������d<M�
����������z�Z����;]�����q[
Oi^ɿ5���K�+]��ôI}�ʓ|P7V�~��}�%�l#�ꊂ@u�#Mk�N�w{��0�D���i��b��f�e����N�i��g�C��8���:x���&|vܶ�f��lS:�#�����6���l2�U<�^'������.Za����ۮf�4BlB'��2s��h�bS�t$�ۚ�;Ng�|�@�� 5ӻԚ�^J����"�Z��0�yݔ˭<��c�!�Gs���DT���	�G8�^�] �����C%v9�=A��Ұ�q_���/w۬�@��x��@H#u�����΃�+B��q�(;i�K}D�G_�S&�_��:K�JQ��d���q@�iCNd�Ar1`@_�)6���sV.Jn�v�b �MO�u9<���Z�#i���+5`�V��Ͼ3�o���y֛^�t����}~��R�#-7����3�Kh���GD罈N��k����ܔ����q�ef�=����(uYR���1��b�.z��8w)˘���=�2�ki��N�y��Q@Ԑ�]�7.'�6Zb}�0���=Z�?N��aáP������ۂ�@�H/�Df��*PSz�a'X<Ɂ��({�����j�vm�#�n#�!�帹�5��WX��b5��H5#C���2l�O��i�!�Y[w������ܧ��1�mdۘ�^u�<WfH����@hGd��t&DD�s_����G�XmZ_�׭b:L��ґ
�1.U􂀁�UH#��ژ3A����0��Q�����?�����X���E��h!�]�W�����GP�mw,�.`�K3khM6X���W�YeIz�e[Q�ܩ`����~ܰ���3n|�nDs.��xX�ː2+gU{"mc�/�s�r�I�^(���,ۍ�?�B��')�?�}��/0Q�z8ϓ ����C�VhNMM��ey�0 ���F��X~[���U��.�k�(�xJxr��2����TD(�&��?��Q'ٕ�ɩhK���O�7��up�{Z�q��!�E In��Mx�uk9�:um{\3��L�2UNhd*�����u0�Уu�=qs�n�{ܭƪW%:-ؐmsx+Q���V��9[{οP� ���w`J�~���~%�����ƈ��Cp  �2vk��������3���"9'���+���X�!�J*�* �<'��(s/�B�w����;q�@�8��"8x�l2	ZQ������m�!=���nʐm�X��lRSJ/���j�ZM_C'*�<�8�����+t>�p����`�<�.�zF��U��ڴ��-o7��_q�>���ߙD�&��j��EnE��YV��JB8�{|�0+�x��Ӎ��i.un��K��dp<�hC�3QDC~V��$���a��q/ѣ"�X3��B�Tl�(9�}�wJ���k���%��ޭ�H����Vfo�����謶����$��x4{+���x�E'EK�J�e� ��A<�j�2C����)~���v����_����Ly�����˩vsEX����.��n�ƨ�u��h�]׫�^�ߦ���'��.�p��l�����P�R��K�:v@�э�Wd���Pb���P0}=�:�5� :T:�1����G�"��ƪ�ኪ���[�K���� ��l1KI����pk�d}}ȍ`B��������x���51KN�6~�4�Jjށ�
6>�³T��8th���{�a���dK!fʓ�4����PJ��}���u�%g%�H�;	��^�@磸�4O� n�9Ħ��\�)�Ͽ$�$h�T)��Sh]?�}`P}ؓQI����:�}ګ���(z�y|����z$B�R�0�e��1�YL-F�:�!�U��zS�2%ru ���h����V;�z��aQT���@av��Kx�H���=&�����I������Zg�^��c�����J%�!����8����וOy��<Ԡ�>WMKFe�c���ڼ F��)��F �T~�+��+����<ʄ.��pk��9>�.O�֣j?�"s/��.��={�C�o��x�������W���Z1�A�94�O��|<_��=q'lf���/�>\�5j�P�j�-�P	n[��M��\�T�ܣ� ����ٜ�� R�u���]ZU�w�$��
}���lG���*�tB��;	��eC;�@���HI�9�S�َ-T�T�a܉����Q-�C�RCPq��&滑@HH�I6���2��-�O��e����T��qd��c�L�=�9������"�'=ĥ�7ks�>v���d�S+FQ�}�k9_��<�hZ��@�*3�*�h�t����ߩӄ�ksv���c�zS����-@�d��aPY!�ҐE���q����n��U=אxA�)�Ew�ó�A
=�|���r!X���o��g�%�º�H�,
�sV�{����|!����`W�_C�3O���P%����>���؄1d��`��읭�!H�Y#��ӥ4�o�ǒ&�6�gqq=*���!�@�������?�i���x)�I���ߧ�Թ����8�-0g�6 h��>��l����?��~C��B3䱻n���`N'��X�B �!��T��=�� &mQb�(w�*�%��Ga"�<�A&$�����)���K`��C.]���$r�Z������p���Α}�q��� ��.=h�}@�"�������A����I��w����J��V��l��	��
���5��ul�j�z�������;�'�=�_��P61�?ϋy���5
5�\k�B��]⩨�����2v./��]X�z��b���v|��Ny�ݴ�4�� �S,]��8�<�o�A֠nV������S�楇���z�\��q��^<�(���s%)g����9))yK	!�8� �l
X�Uqw��	ˑ�|	��Vs��`�[�b���Z�/��!Hc
���;�ʿR����Lkq"{ն3z$g	}�u�[�jfG Qܭ��;���>h�}��ޒ܁�޵o������~p{�~R�8N�i� gp�;g�)Ӻ@u}��{Ag3mڟ0��z��y�@0�hrx�����,�oq��*gp����e����RF��钔�U~"��ᗺB�y\��7�*l�+�Z,��qY�
�*�3Ȫ��o��ʠ팃�N��^�����2j#��U� �=��=�a������H�v�a!Qy�?�La!����;f�ռ|i�*����bh�e��t�Lz����Y"e�KG���x��?���6BH?�[�(�#c+=v��}�ntoaj,O�e���I�����Lb���ͨ܋�6��/p�V+��[��)��!Ї\�i���[�@��88��%�{�hE4�*.F��%�N� �f'�HTl���d�F-�NT0�pT���m��,,���j�>U �7��̵���"EY�_����ᲈe<�
�$��`�R��F	ՉRgcw�-�Ap<2+��ok�hjj�Q���w�i��r�,�Z?J��q�Xs~�O�;]c�'/�6\��-��YyFF.��;��tsʶ�`b��2�ȝ��Q��x�ޣ�*Zj3�϶)���?DO�,�q.���(��vc0�w��\5�V��}�����
����Nz��ȡ% _k���"��?%u�� ��=3�:��$���Ƭt��K�:�sM�I�h�B8>��W�.�|�5p���5k�7�8�(�k���s(�l�#j�����#�!��̿Q��)Ǉ�{�?� �h��v���\u�������0�C��Om���� \B�{q�**�6萑��J�R�tb�٨Ry�*;�E�H���;�+�Ɤ�q����)�O��<�	�&6� ��H��u<�7w�ױ�x�}���Y��-!��t��
z'Vs�c����^�Z�ڵRi��Q��6��;�{���k"`<Lw��"��k��TR9�7=��@u��҄ylȧ��VI���~���)���/�?e��Ј�e��)$�Ie��i*hh~��S�',�]�o d��:>�5�X�7��A9_�K������qt�Ix�c�������Y��@�On�E�G��mu,+�ð��E�N��!�#LV�*ʀ��;�(��%��]jt䮜5u�<��_+0�k����˯��%Y�q}eڒ��h��>�o�_�^���ׂ@���=�I4��'�Q��ڌ�����9�)34�z�@�$K�|<�����7'qI�;!� pރ7�j�$��N�>E�����6�tZ@ц�i�"�+M���N�l�^��?�9j6�N�@���e3d���<�H��qHu^Ñ�3���H�z�����k�IA�q��Ϫ ��f�x�I�t3׾1�g'E���W�����M><QE�w�F�X�'r��g��@!f�d}�l�x����^6P�� 'c.��>����!!�
%�h�bgr��ސbd���|�!|'pK��)�+�/�D�|A�&.�8�I�������ҏ<L����j�l��o}��.*tE�l,��ml��,b3(����C�	����Q̕��ᔏI�W���@��� �EXtŹ�pS��Je��1�Nw(�z��n�4�XON���ﲹו�0���F��w����/R�)��,����8�B,�;�5,3-��c��ҭ������:Օja�Ex*�D��n��������m_��0���Ӵ�Qx�������?�x�7Q�r�ѵR�M����J��s!�	�`�v�``�K�׃���;�8
�>(��r� ���l��|`m3�����^A��h:d��P�4�9rD1�]�A��l���^Md�+�_�6a}X�����
�T2�ff����>�������[�@����Жd���j�g/��Q��ְSx���*����5J�6�yO�����@� M�a$8��>�L��:<~p�|�!,�D�t��*��/|C|D�ҝ�8T��	1Ȋ���)�����H�p��p�����M }�9ȳq�4f����Pb5����YGu6��j��_��wс��v}�A �'/d;*��zZ�혁78��+H��a ���7�8"�i��֨��~�&,d&��i�>�Z�Ì/�E���0Y��C"����,&�v��ֶ��N�9���N&��B�o��e�3��j�n�kJc�<��4g����I����,�l����ai�˭崲y��qB6�_?{_u޵���;�f�7�g�>���6�Y!$�a��)���C���Q�P��-e��*���nx-�wOj�:@�
�l`jAnN�"���ڹ'�<ͥh�v�qc��F�tU�] ��������c�F6��r�pH�L ��
쟆��K��3�̪�D={`0�"<qc#�Yf�"Ǖ�`�$�D�!�h����4�� ͡�Ν�sL1g]pCbYO��I�$�/���2t��:�3>Z��_��:�#�)�\��P�걀��x�	��P�?r@��OV�/�?
���e�� 7(mC[|� �Lܩ`����ޢ`x��M�� ���x ,&nEީ<�;6y�Jа<��4���-��	������Q��2���XZ�C�}Z��70^�g�q=��6���Ŕ�����g_�[ ��E��B�a���c�WɃ�^�@�8f������]� �6�Ǯ��=W��0"�EZ��q!�쬕����E|�$�X+(Wr�;�����6b��p\�-���i�ˑ�z�k���)mW��덪,�b�=��$ݚ�g�	w�w���F�|Z���v��X�=�!"goO�VѐF��V:���� Q���y��H��'��^m6٘���ۧ��j���rS���ZG�(Ld�a��ų�y��]�Zؠ�ĵx���̪iw�Sn�������+�tʕ�QE�߆��>5�J{Q��^W��>�M%�1�����vRn���%x]���3ny������.�v�_ˎJEE$w֏}�?|U�s��Aa{�}3�|9(�i��輔{����u�,3��au��0��bF�#�V
*po�wu"����d��:2�,,���^WPa����r�d�^m���#-�g�����&r�#�a�ee�� ����߂"ڛ&��[ƚ%c��%��UP�TS�m�������졪ц��A��EG�7��6h�"��28�g��c�P��8?���V���*B��-*p�Nή�g���e�&��l�����*���FZw>@������?�?L�եXH|�cN~ֹB�D���Q��Y�����)�w$�<��뫫��Z��,�/�D�+��,�GA*�	JG%�0�YX�KOM�Da:�x@���%���ѷ2�Ob�pBx�Љ�<��	�
B�T �E+�m�4��7�jҠ�d"H����_0;:yf�{�-^�;Jn��77u܍$�#<!Z��O� a<�$�u�̩�6�6 Ď�tۮ#�faH�J(Po$:�H~bT�u���KW�
i�!+�D���_�h&|&k��Y�M�+�X��n�x[�u��3�ݵH���v.W^5{�+	�U�{��_ŜW��V�SSB:3�~(be`��͖���l��h��h��m�K	��Q�O`���b�P��`q�Z=Ny��~5	�G㍑�F��-Ƀ�ͻ�YF���0G2�^!��ɖ���q_���Ha����5Q;6y �Խ���^/m�8�y���$#y�Dd�jRfH]\-�x�c~�/\X�K����DT�D���U�$(�]�*�<.��FL�T����}�����r��F.8�h�������`��7���<��� P��f�WhZT�D��+5{*�'�$�H�/\=�2A��S�u�U�ǒ�U���d 6���r1��I�כ�;SN2��&26�Rm��jʚ�K�!A�lh�~�{8�>5Nڠ���5���?��_��'��1p;iW�+~�i2�vٮ��i�"1��6	��x6��0}{���g�����'.35�!g����d����L�J��*yK�d�`"H�]�Q����L���]�6Ģ��� �7:>54wMq=���B'V���o�����`�ƓDX,�ȋ�m7� t�U��\YN-�t^�nv�ܨ8�U8��_�8�op�ٗU�� �3$":�7����M`����T0��X�@-�E���j���Q��������k�# ��nyeU�2�N�Hp����Y��ܑ�;�a���� ,�z�9�_j�bWKC���	L�hF�ki�f�
����"`&�b�b����hbR�$IF(Йr��0�y�'��G��u��+Cg@deV����[B#P��Qh@��l>�J�����P�]GU��}!,g(+��"�4�%ry�xv���5��W���8B�#DG󒔆c�cH:?�D���3�My��˱=�h$��m��r��5�ŗ��H$��m�:���t
񰩤���Sq0�x
��ü_dDlN:W$�d�n|��Nܳ��ض�Q����S�oqz�A��c!ؓT�60]|�6e���Y(����2>p��S�4V� �<Kv����$)Ċ �
/ș��y8�Mmz��׊�Y0�Ô�� �74ٶ&AQAA|͚-i��oVz��&I�}���ZK���=C���u��0#����ӌ��۲0���d�ͥ̂�%KzZ~��u)�w�"��/SQR�4;<�FLʞ~h�\�'(ReF\���m��ud;���Gs���kUD�j��	V��'�؂
�׷�ހ䏍*� m�sa?0¼y�:��	���ފ�eK3�S�Ң3�nV�V
	i�ځ�E�Q�j	q	7ݣb>�er�I�.�g�c ���ᡸetШտ{$�O�~���w�;�;��\���ռ�}�OBf����4/��c$���>s��FT�70��9��$(1�mur6�Qzj�ֿkW�I�N8� j��r����1�c�s��h� }3�2�lG���[�:����{�(Lϧ���e�>��c�����@��X$���v�VE���6���Tk.�՛���²����n�:����i�l2}��T�[1SV��j��]�8'�y�[<}mI%���k���P�&O���ZΌE�����ʒ$�)��k���8[`x��hշ𢹷H4��D瞗H���)Ӏ|0,�|���q��O��nXC����sj���;�s{&�S����̾��8�"'��
/������4c���"���W��%D��L���jSTQJ�ǥ$T�p�	1��۪�ޑ,QL�(H������nӲptV�+0��7tMMm�>T)ʯ[�]a���AӲ:P���)������W63YZ�i��PC�T
է�I��!^^��~B���i����whkў�G��`�B,� 8��8^���فu�I�����-웜��� #S-����;:�2� ����"��Z��#;�E����v�gC %�SfM�p�;�.�WZŜ�C����=w�
��PE��O���o��=��A�;Pb�ЂǙ�+uF	�VE
�f�W��٢V�q�-��ʦ���^���?̹rwe�g1�R#��̿v���1�W�YM�?�������J�ӕ/�4#���W�`�^��i%��G��b�Aqx�7�M@|�%���t>}�C�@B��Ç�qfb
D�0Ƀ� �Qa�,�e�?�&K�,��������dǞ��O�wp�SV8s��:�f��� �ܓD��Ɋ�n�i?�?|0��@Ӱ��|������A`�9XFm�g\zV77� '�r�߲U�s�Z��4n"S�sw���D?�/�'i%�4sŤhu�ξ=���U޴(����CAa�Fݦ]1Q�t;��G0R�ٕ@Z�n;M�-V��@���U�G	��S��>_�o�r��j�!�DP]=K��E[���b����cI�hL�L�4��މj8�&��4!y3xs
��o�����{LWb�x���sFS�/�t^�?O�V=�٠@CiI�آ�����֋g�x4�r֘W9�<a�mh_�T%�v# oP�	���~=뜩��5�����Z�Ks����w��G�ۙ�]�bM��*v:�}&����2��]�r��8R@F�~�|�漲��!;��]RZ�y�G�Mqf)�Nk1EY�*�z��6]�
����'� �J��⨘as	�=/�jݓ\����h�]�����K�sG�����4O�ʂ�%�}�ʼր����&��I�"�=K��Ru���MO��ƶi��.4|�H�S�!�1�,�T��+��Cf�DG>�]�����DUUm/8W;�N����}��d@"@Ym) �DE�T�A��띨�����"E<0ފ�煐�?�6��y!���+]
m��g<�hF�ǻ�#���]���@�vZu���j\m+m�� D#��h釻_��Kk�x�w_�������^���E9�DL��Zɛ�KN�|��J9�c��$���f����� ԓ.��H?P=�j��t���a�䖪m?b^��:b��A.o N�������l�|���K=HVc��^�y\�Y����da�$u|`��@��E"��^�颒W7QmC�d��~�������I�h��jd[�C]�t�*BA6��z7��'<�H���c�y�8��꿤�3�p��sT�C6*_o2c�M�_�P&���x2���S��q�_��;��Rj�㝾Ġ��ӁԪ3#5���H�&��� �eM���cs�*=0^�sR�,l�;�&Fx�<=��#.:[��ق��x�+�-�n���P X`D�QP�������5�|.0z1����Ŧ9�t��n�%n(k�Ug*�p�Ш��G�,��Wfא���'�Y�89`z�����;t�J4!�_~Wt�تQͤ�+�?b��0��)���fz�������dt�pHP�A��ڞ��y�C��_R��X�:ʣ��
_�+$\�"�(!���\��R�OxkB`�jn��N���S}�x���XtV�����+V릐K�9�S���:8_�R4m���o8h{zb�O��x�A�+���R��]�� *�<�sg����w�Z���a�(�Y(�Q�.�;:4A%�[6}ڬah�M��1]ԫ�{���#o�}�U#��<���E��7�%D����4r������e��	�O�>���v�}9���WV`nR���Ƀ9�d!��"��S���,���l[�~�����F ���t��#�i����6�ӵJ>)�krq�6x�E��41�	\(p/TlT�s<�p�M�y���5�h��uL7h�B�����i��'�?���ԟY�"<ǽ���Nf�舟�[;�~nr%���òM�3J&�3BRΚ��"1�$��) ��K����˰i\���6��Q�'�9�?q{�k��Ѭޛ@+P(ɦQzY o�S����s5K�d��}`5��Ƞl
X}W�t��,�U�z ���m�E�����c�xsh�U]�Ǭ�踡���?kҫ\��"C�C����~&�S-�jSo3�)v����T7���J1.�Y�GτN�p�
Y&�[U�;f_�
�ߚV�*��S���%�j��՞.1͝��У��1�c}�����|Ԥ4��e) P�f��?����n�,�1�,+~�_d����n��@}fu�}..��N�4�����/���PJ_�T��Gɠ�w�!Ke4l�ch���0V��P�U�;&� i��3Mb��}�E���m,��ڡ������곅(��&_H��*�����N;�+.2��!񢖁I���y�|�KN3���y~�_l厇7�����"�z�6���'�a�^����ӌ����oP�����?�9�y�M��,��.y~P�Kh�z���f?��J��2J[u��gil'�Er\��1�7���WϏ���[&>��(��7Y�7�ߝZ�\��%�WJ��~ԟ�����Ӓ��l,���.b� ��tܣb���Y�����>���id���Kru��x�	���N�Lc�VV�x
�@\q�ے[����k��>E?bd��+W2A�ȯtf@�f�N*���>�B��i�a��F�^��5"��)>��F|�&Υ+%m�,i���a��]�z{�͵��K] �"f�~+�vPW�ߥ�z@�Xi��j�v�g.��Y�ǣֶK3���Dwxf[����(�P�mD��C~kz�� uJ�����ݝ�/`/P�}�jZ<7�Qo��B��&@bo<���tH������.���2V% e���<���9�����[W3՝!�B��P�y�ϋÌ(�l�ڎ���1*f�睝�ۛac�0F�bW�L��&N'��4ڙ�=��W���VQ�[5��K�ǯX�]3�wZ�{�M'�h��U�&%�SC�o�'��y3'�s��9� (���4�����K��u�����_���qJ�ӁI�j$�͘@ W��}�mۏ=)L��#�v8:_�����[>���+�a�ۊ\̜��^�죿��^Sq�c���ukt��9���Ja;�3}��5u�Oѓ�籏�a.MTX�s�%���(��쓁��}�gx����V��t��Mk�WT\��s����E>9�,����(z��o^��] ��Cة��'��S��wB�/ރ�ɘf�e�m<s����\�rof����UD��}B�׈e9���T��_�g�Kpx���J<N��8��t�3��;@�3c��|�s�<^��GU)�ð`�D��.frKZQ�s��>�ZS�iuI}����TM�){˶���;L�xه\�)<d�S���D1w>�tI9Q�s�"��HZ��4�
"Hm^zpu�� �u(�V���5�%-����xZ�*��H�e�`?]<�'�e�k�Eף${,R�h�"Nt�F�OVg�`5���μ�rQ^�^��.b�f媻m����F4�'����%��Nw��N�4�A��<J&'�z�cӴ
`9�)5X���N�eUR��Ռ��P'�n��?��"O�.T�
޶
��K�Mb�M��E��k�	x�"X�_�%��m~L����;	p�K�WV��;l��/9�,r�r�$ӷ=6N��:N�$�q$l3��g�lڃ���δcXw	��|���ٗ�+Db�4�b\Z��ʡ{X���BY��c�T�O��R��I-lV���ڑ}�%�	8�5h�R���U2th�i6vB�A����� m,ӒJ�t��`��P'��+I�F����W�$�7�o���u�뱊��`}��\����$K�a̰�'�-���L��yڻ�-��k�,!�#|3r�[U��p���� ��G!�"�4Ʈ}���|}bJ���]1���$�V~}��E&%xэ�.'<Ψ�LF)�� xTXT�Os� ��Gm��� :�#�vS�Ⰰ :�����ާ(q��ks�Q��\YA#'3�ܥ��De����PU��
:t�|d��l3ZP�%�_9�k�kӢl��ȹe�"�
�s�;�H�_@tz���z@hOr�&�������.&�/������3�F��:
��Y�Tj�ۚ���6Cs���w^�2�]�b���p�X�Glr�cJj��Ib:3�Vf�3�5)������[[�%�O�xP�_O�v�1=m��#�[��v�ߍ�1�xx�^��F�������C��Inع���+�D�49�kύls����N�?��8�b���V[�`�f�~U9q�	�gm&Jyw���S1��I6B@ql�ӷƍ��;v�b;�&>+�ԗ׬SSӸ�u��[�'wZ�~��C纵�{l��&e�iM7րqCȂO��9�l��v T��$}�?ꝩ��*�&��yz��-I�u�<�@�u�p� ��Nk������BT�9)���39�!�N}��)��p��?L!��� �~E����ULrS�*%�[�����d-W�� �s�JG�i�qV�tw�&�3"�eAW���s� �f� ���k���*~UMk�F8��+�8�6��,!!ӓB	��`^�`�)m����u�IGS�"�d0��hK��E����y����j[�Z�}��@�|�����(�`W&��b�Z�����N�̀�9�n�a�G2�<"ȯ�`8�A�R�=F�ɿ8*���}���q�?�tQ�v�0��egB�_�.�E�=��Nt��o����`̧��b�?�6��l��&.�{����P�ŎIe������ާ�h5�ک��i$��9S�uY�Y��%�Ǌ���q���k��S[B�|�]�:9Ks�����
���E}T�1c���|W/�]Y���MɆ�uu!���ͮ�m��=Q����Y�5|���ǟ�%[Y�!J��v��謹xRPL/Ձ���gEn�`R���JF"��%����&i�!��s�e��So���
�I8�Ȩ.����
��|���G���&�����hӝ]\�3��
&h�	bK�D�$����	����ǙGוqd�c�w�K!⚞���~y���g�C��u�8�Z1E<���^C/Q{�'�t�nT���G��Y�B��N]�υr�x
���ٿ��:8�;uf4�z���<�ǉ�<�(glf�oΘ�*T�X�9 �6�`j9I'��#��H(�G����!�Zt����7��牔�6�w�ԣ�`�z�.��'������u+�=����a2U ��'�^���H.���y��9��o^��h�i���-����3p�ZL2�r�J/�|q-��_���E(������U*Ӡ��4��]���u��%f {�6�D���td!�7�Y�;u+��'س�f�Iq{�(U�E�UE�Y;�\�2HxHZ�+��k��\�5�gU����aln�h1�1�Q����k��1�.ɵ�}n���|�3LD��+�)�q6��|���{�2F�|@6�`���
���i�������$��-�U�`�|4Uao��X���(��P�=H�N�l�c[Xl^�}is{	6krk�WC4���soo��fT���-�<����MN�~���8!�R\�A�td�����o�lŅ��?Zl	�>b���G9*K�~�+�a��XH��8/�|_��8Ԡ�F�K�v��M��OnƋ-�e��twTv��&[��H_EJ]���{%�P�%�/S��2���^����އ�N��kA��E�:3������>.�N��q8x�_yI̋hmu.�]i"}�SG%�f��f�����8�-�����ЕqI���g��c��A�ۥ>zT�8�K*L�~���$�B�����v+K*$G���RSa������������/2���;�+��y7c��Kb�����,�0�QL߻G�mv+�|�چ<h	����ɍ����Y�x+J�_;8�Xg�*m*]'|o��Λ��rq9�Gg�'!��@+-����Q`��EL��qԜ���S7d�rY����<��R2�G�yHF�0�|�ʱ��a�(<�+u����vM;'�p�pS���D۽V�H�ϔ��."C�����t�f�h�tt��8�'�IV�,�G��ȔΉa�r���2<��q�mb�tt0�� `N(Iں���>�-SPč/�=M�����g�J�,!���0�w,���� 6_F	�����Yfr��v��о1<l���]u�۸�σVq\e�W�Ķ����~��O�r��զq��E%�C�Ѝ�+�?��4�rRY�9ل7tY��� ��,!d�5�@�6��Bz�;�2[K�q��X/�.K�6j��9��3f�lr�>�3�oV�HS:Q�`��˱6���^KB0��=+9�Y�C�iS2Н9�D4�5�b!�d��{=e%d��{U���%�-zs��SF�d6���i��M�.L��s��ǉ���g�:�H���Ȕ���6�)|>T7�gE��__�@�l���$��
����3��yP.��%R�ME%�<_1�Kq-�RZ������Z�*�E���c$\m鞒h[�gP�����"�
�U"Ќ�,8׊C�s�朽c�)���?��ު�p�tpO��tG˻��jTaU䄍le\ 9<�_��<��c�z�r%2�@:��cC� �T�ig?���K���U?
�b�γ�Qc>�>DV��#��^��i2m���wv=G��qF�����< �7~���d�'<��ýqg�>~��~����@�
����R�{�H�7��-���ɤt֕=�T	F��b�u�H۞������'J�v��{pVz�7�єS����@ �N�UDe���sE� ӽ��Y_]_٥3v4kߝb���<`k��r�S�Qs9]6P�=a�:���c�)
�h}��qz k�
��]Ƙ_tJ�w�߅Qk@u���k����k��8�&b7w}��F�D�h�xf�j�PN�,���������z�:�н<��>x1����Կ�)�����4Oq�Z�=P ȼ_����c�f�=i�j���te��aڦ\����F#̆2r-��X�����O��2c(���	+^�~9m_����',�`@D��OP�d7י��/)�j�U��E'M��q�e�����U�.� r���UZH��(��Y����"���P%x#��-Ќ\��h6�QY&@���:�)����F�S�6����J��.�;}��`�h��`����L�:�$���w/�p;��(�m��������_VgCQ����<�v=^5e�4���V��� ~ʲE-_Z�i���Yn�˹�D1���F��˩o���C/N��g��an�b�����w3|�R�{����eh��WHZ/'���ʫ6�<�w�#@H/q%~>�����B��ze��KMok�͉�~���H�����<L�U'v���fS�0(�$j�u��~��Y|�"o���u0�h.��	���o��XU]5�;.�W�·:t���yy��UY��v��b�A�C��	���U����N�rqksfC�+�����6*�����n{�}��JoQ��܆�-_Bf*������$�F�m��+m��(Hф��D������gn�)��{���6W6��a�!�0@���t�it�
�n�\{z��L�L�x�m���0z��<}8�u�P"��U��ao�=����$��J�<P�b��Q�[4*��2�g�gv��Fv�[�b�Pl�BQ ����^��}+�3�{󷝬����h�t��ۈd��{�� .\�̄�"x`[��jH�=��%P�8Q���@-�$ ��4�=D�N�eԊ��?'r�4Dk���ܕyH��'CB"6�;I�*��17�t�Q!l��KG:V�T��|�Ϝd\rV�
��=f�[h�}K��lN���;�_^�^Y8�S-��Rl����,�pFE��F{(J�E![���>8v��}^>g4�9��a�|�Ȅ��%����{�bz�1&�V�!��q��eM8�\ �O꾦�.*���˽�e�z��gdY�*:�Ul�pbQ�qXڒ� %��|�QGV���>qv�b}�8#$Q�Y\{�֝t���*�uUn�=��#�p�#�*w`�zDf�l���[�%e,)�9זFn���%cG�KE�U���o�"����=��E�nJ���G��7����M���W�Z��"M	��w�o���>q!��w�>$���PD�j�t'X����g�#�??>��D�EF@[�x��KY��?���=��'EY�QG1���R�5?6���O��a���.Tn�zq�}&�Ik5ā
).��oƗ�AsH���N��h�e�(�U#�.�ٹ/j��q+�^%%������d|��[Ca1���4Z��o�]*!�>������H���lw�|�)4٧2���`�B%�ƿ�G 7�����������I�ƠPHh7�*0�*�F	�u-W�)a�����s�����Q1H��W>���8��>�5�]��']5VZx�ɧz��J��S�b�.�y&^X|�DB���7�vA� �V:"
�l��w��C�;��V)8_lĬu�::���0I��د����TRد�+G�d]�K�C��7C�j�u�4���;�9��	�0�ë��d35~��4IM9�"1���_N3B�y��m-��F��=�Rl�uPĔr�^r�#�s7.|BИ�k���`v5,Q�V�jt�/����[���c2�v�u<	>�i4��L��3ߠ��@��P7�#A���;nw�"���	l)�=�,6&M�&C�I��n�<dQ����eP�Tar��� ��1��/���t���Q�0��@�$|��Hc1�}$����P'�"��+.߇<@z����~=0��C�E��78fEuA��y��KY�C��3����xF���O�p��\~�/��[sa�~��?�iW�F.���Bv'O�i>]�&��9#^B/s?��9�:
ݖ���t�\��8�<vO����<���?n�̬v��/E?�4-O���l����	�*�n�b
I,�n�������2��q��a���P���sc�\a�4�N5��}lpN����{l�9 ��
�I]�F�r��c�)Kk����=ؾw���}���~HY�7)�4ϡe��q:�l�z�����|��t�-�.� ��o�����0z�ݻ����=���nNj��[p7� ͕�_K{u���"�]Ep~�{�W�H�����QΈ���ï����nx��l|��@Y�j����'�����z�m��7�#�~o�-��e<E	 I�p�-�L���2(�fN�Y�V�Mp����eeS�Vج�m8mW��Wg���u�%fTw�҅�7�W�Xv��ԥQN�z1����/��t�����zF�-h��5�2(T`����h��,��Zi;uiN��9)����:�
t͆�kE���Ns�}&���O�3�!�4(!�92��[=�!��qŠ��kۡ�XV�TR��t�<���!<{lᔪ�)N^�^U��m1�4侑3��5@a�lic�T�
F|2	Fz$8`ե	�lg����<A~�f�)�)O��+�a�@�)W/��xϱ���}汮4��)��^���ļr A�z2t�Ȁ5R_kd<+�e�2���D6[�XJPZ���6��5��'��-·���1��c�1�ow^�&��ib [����&h��U��y-`��oT���aO������ny���U�Kǳa��ƈN�Pu��Y��y0>�s!���@+ߊJŶ�'�A�W4�͝���]����0K��O�qɪ��p��ɛsM�9��鋤C&��r�r|���i|�$�[Q~��'���p���,n��z���B�M�V�b/[ݭ��ԛ�'�ˇQ������� <�p�;�N���K!:A�����%k9{`�o�_\e������N��`X2��4L��fa��ӱ^ :�w^dp��|Ϳm� �+���_�;���Y;1.qTmB*�n�bM�,-)��U}\t,�՜��5^߿Ӫ�y���u��`ߞ6O�MYvG�f�\�D���O�q./�ciBJS��V.Ƌ�qC6_��Zk{GQ'Ko���,ƭSTk�In؇�m �yז��^)	����^�YEA�����_�݀c?�i��!#��T���%�[�vl_aE�B6f�[d.�ݹ;S(�
!襶����[�]2"�~�<�QLQ�3ޟ"����Wd4D��?x+e��a��t�\=ʉ�j��'�5"�Ƃwǵ��Us����<�џ>6�i��55��l<��'�r�T� �I�u`�m�絘� �;ޜ9��ORd̍�� ���t��`5�{6���Kw�� >4!$�g�e.>��ժb�#�eЕ��!�:M�b-l�J���D>�meh�x����r5�O�B����8r*Z�a��T;m0���J�W*��γ�֔���Q���ʀ�c�_��L :��ۢ�n]X���H���u��j(���2��$�XgcZ/�Rg�	��R���8�� <�Z0�(�<�</�o�|�j�L����e��c��c^΀[JԞR֡@38YCT�dv��f~�gE�0TX��z��?�zPCIA�9N����L�*��h��1��+h���M�J��Sz�p�[+���
�̝!�n�}E;���BE��1���jo&�����U��L]� �v�ֺǿ"O��.�m#~L2�,�����-��:�:w��.)l'�.B/.�0�+�}���:-���h�w��ܑ�)%�L#$	�9ѭ�PR�kj��8��R�X�H}_V1[ӊ��!�5"t��H��<�5Kt��׽n��/P4�R|SMt6<Z���KL�mc ��w�����s��g�`4/L�`1�>�B��t� ��M	�|~�U������L������_E������Ǿ��s�/+M?��&��_��Q,ep[!����֤�e�H��x��IYX;WW��8�h2�]�6�Y�酌Pp^���疭6SFsT.�ёB���3i3�����Fd���/�$;W��(����!q�s���n�A��cAx��u�0�NOa�{�����j��!�uY%��sR��*ԯ�����
&�H���VY���ǵM�V��{���}u���'	�_����`�̗}̪<t�=�n@mm�J�ڼ�ؠ2�^z�`�����Z�ua,��-��@��ɒW٥aE�5~���`�}�r�O�����O�8A�e���&� ��Š����Dd�1����'�mӺyϨ(�
�@uby
���������dO?�,��"�&훕5kТ��T�Bm1�5��A���� ���/T||�;Y�eS��}G?AB۲�吸�E�~N[Aw��0�R�0Ę�ލ�%����܉�$��an�5�&*���X
�^��:H��ҷ�Y ��"�ZJ�UpGR�Bf[|���$φ�t�����q��^+�ҬfLh��p;��4i ^����@�>�-�F�e���,��5|C꪿�RxݺUyO�;�,�ΙZ U�,[g7��
a*�ھ�kH�]���bxŵ������ϩ���p6�x�+<'&@���@/ �ѳ�e8�Hq ��"B\F�f�L��۱����h�?F��م�+�96�Nkj�S)B��/��[D��;e�VU��Q��Ծ�ܟ��<J�n��ԉV��,�*��ο�j�\�K4�zA�f���q�^��cZ��}fdeJh�A���n�y �?�]�����������c�n�F ���R�%x��"6��9��nF_��U����`��RoE]�^���b����I��:�킔�╙Q�n�`����:z��2w�;�A��l�&_b���DsĂ��+L�@��/�k]>yi�ZW��}�h��;Q�%�|�x�]�����=}X� ����ak�Ոiv*C��Y����{�(1ǯ�l�3�~�H��x?�g^iz&�=�.�e�]���-r��ybh��_z� ��X�B��k~[H]]��:��=�L�:���h+��\mj6�y��|1��}+j��J�3��+7nS$z�s���'��alT��5��̷^%�vr݄`D�:
�`:ƺ �o���B���{ߒ�Ep}e����ط8��d�(V�6��cH2��Ǟ���C�g�$�_l*04�/���	 =@gcƟ���wqk1�-��{�%�"yS�z������vVT3R��>0Jb0q�PLS6,]��4_�9��u���G�^�-S�po������@:ٱ�Z�S~U3��t�,a߅�.b앍���:0�����Q�}۰Ni�l���|}�h_.�2��#�S�=g*�.ֺe
�(dsT?	O{1�ӯ~=0��R��!�I�-	�3۫�҃Y���8m��*G���ε����dk�ͶUg)�iZ��b ��.D)=��sH������^�[�s)�6����)�σ�t��
�I����ɰv0����:|2�!�LV޳���f�=�1�'Lz�dg���C6ٛ�IH���w3݆y1H�"�!o�s����)�%t�K��ӂ��O�؇@�d:]u��	Bv��|6x1����(r�o� ��r���yAflǔx�Զ��LR�?3'��5�[U̚2����1�N�����p�`nZ5���v,����V�L��(Gd
��8P��q�@rc���9�	���"N����;�`�B�b|��=<��� ��a7y<^���!]W7�o�D�0W�&&�Vh;�1���4"p��ҌѪ���]�� SK��Wls�[�JgX���O�Tl5��F"k�s�L�2B�Z�O��(��l���}������S1�Ԭ������o���um�[.�Ƌt,�!*ڲ|�L#��2��j�����أ��x0�%�ZD�-b�m<�(���������q�>  ��B��&��v�@������}&������8�%�kŤ�<"�r�w6=I�� ����k(�a���U��Hm���I��@��z3�A��1��HU�)�Fh*���5BM�i��>C�Y�m��p1pJ��"6fl,.�#�y��:)'�WF��N�I��wo�����*P�.�.���.^7T�P���J[�ST!K���� ��� 7����{681���ל��7
ՌAB�_j�����7V�ޟ����D��P�u]k����ڿ,��R����R�!���S��]sٰ0H�3� N����_��Y�Nķ�k"6O����u��~X��q�D�a"��r�à��ᔂBʻ�A �l��&��0��$��:�ѺQ8< ��Aw����Z6���lF~J��S�(�Vn�]��+rd|�5��䏏�S�q���On��2�C�T%�,���Ay�R�wK��{��3���s�c���6���$�a�Bq������9���:�p"���	z1��CXk{E)_B�j�7��+�W�
�>]��*<�����#n�����DKkQ��!�vg..�T�R���AT��D�Xf�+��h��E�Kڰ� {�ñ/�(c��E��6�O�g:=٢�;z�o`����9h�[�!�p���B�_�>c_���g0��R_�4��|dl�|�=����'0p@�˒\^��KV���9rg�K7V�k�6�Y���i��\�� ^eH�-_7�#>7Riq�W
`���w�?��msT	$O����ց-z��k�y��,��j�q:H���E]Y{�kB,n�W����]�ky����R*�n8��2��1�?
��v�<=����hB��=�|¦?�
7�pr�bU�"�y����H�8]���]�Z�E��Ɔ{m������j��e|�-����ӣ.�X��K��S��X�T�J\OF�O�zO���~�����_�v_F8\<���XA�&�/	Y�����(fOt[�����Yje����H����{_A=�"�=���c5F-�3"@�ų���Շ&�5i���X�@�I�;7_*ٹ"��JRڼ]�ը�P�>��3���<�=��j�A��'�-���C��[�r>�Ӿ�3�ym�u���L�˻�=&I�v�b@J9�9��U���	����2�\H�*��Ncs��������t3. �
!x����:�"D���(?h�#��s��nh���������9�A���L׬��ɵ����X�.q�~]C��p뛴�$NU�&��p��&#�X�/TIp����魶`�V�k�B�g�CcȧQ��M�q��1�V2݋)A����L����m����5�M�`�o�T��
/�ڃx�b�������n#�3��Jl�Mc4��)�}�ܪ�i�i���������RI��)NZ�w�v�i��<�H&���]��.�'�$�*�Z�z��	L[��RLH"�൤��7�o4��q�.h�;�w��#}[�{��Y=P*�VS&��A�It���ٳ����XR:�K�,�,=`8��F8N�P�U�$��_յ"�
��-���{Q\RYhq��43`�W!��2���5��YјGM�_Ȣo\�_t���RB:įp��(5~t��n�r���ͺ�;�+N�\��{۾YX���Lx!Ħ��T��3u8�+"������ڣ��Q���ʧ�� �V߸�}G_����3"�&��>��%%�%�nH<U�V�T1s5m�`B@d�;'#���/+RC��E�yE���������� N�^@}��Ou�IhU���yՀv�
=���l����!��O�!q���M�*��h��ZRG��(y�.2QF�o��!����@���M�QUgvʫ�@��佦I�/mQd���h��^>��'�@el�V�v��I9N َ3�Oi?��c�*H0129~r.(�����3!`���a&�Pءfgҏ7�>���.j�6�hMw q̓�7�G�[AX#Q7��: �Gdef��y�H ���$#ǫ*B\L�PЮYh2�MzW"`q��[�Js��pRe����%�[_�e��:Yߑ{��{ѷ�T߷th#l̺p��s�mh9�`���g��i��K����Wc���/
��d�=j>f��$QkI[&DF"9e�1�4Ul�9ۺ( 9~:dY<b�q|�*e�i�2��)�,�/W8Ԣ��*N#D@T�vi{2R����g�H��������#_�6(�W�a�y�qЛJ؟~�9:�k^�:���IX�P�]�������JZXL����+|9FG�R-��Tl f济��<��s7>N��f�a.A�W�&#p֧0�/-z�x��S{�#6�EI�D_?���-�*	����kb���b>����AC6���v�Ë
zD�#�ߛ��W�	����Qs�
���s���ѥԦ�N �E�(�b�DS[��R�25�uIx醊?�,�vg	�Vf�0n���S�1�b�]#K�X��$Y����_�E�d�[%��1 =�M ����L��h�)�v�趺��:�x�s#�CM��E�*e�B�ў���%����z�2����?�d  ��y�g��}��E�'D�';d�&i"��})��.4�\"�k0�D�E�O��0酥v:���#�1A�p��D�����Pƚ��t��U -]'	PэZ��功���j�� �^an �ɓ��	�/��w/����@�����n���,��ћ���-s��3��5Rj�?H��Q�)iA-ğ�@���E��`�c�����%���̜�E�.��:��t�"^+��
>K6�mܠ��p���
E�6S�a��	���@xF.�v�C�,�0P�����&ҷ���q�\���,�sY��d�+�YԆ:d�Y�C�	���jj�@ϥuމ��?lݥ�n�{^��?�偔`���W<1�� Gv!������.M?��U����u� '���(W:W��w�r��2�`i0��͙���D��,럎%��Q�w�[�+r&��M�/u
���1�d��~҄@��c����S��a���w/K����2��[�fa������d7J�
��M��C1:0��^���2{�/���w�}�������%����ns[_qy�*/��*�E�m�P(�q�����Roc�_oS��x�5j����B�&�VB	U���S���(��{@�L�$��3#�� w�@E���ڏ=ĸ`*��z���L�x@�*�̛کSH�W���w����]�U+���D�o���wdr�_$�4�������������o�MV9[D�:�!��������I���.<Dc����|U��R�+W������%�t�8Xp����.�㩑�u���n�.j�QY�������J4�_��!�s���1�5p�	��L�r;����fq�f�#y�O�j�X�e�⡅Y`��=���q�Dd)�4���d
62��>P��S�h��!|A�Z�N	��Q�C��,�c����	~��Y�g#U��sF��S��,��H�,�����k��Z��"/�O��4b˚e�=U�AQH�M���/�Q�zq�j��-���I<�4�mdg���q�����4���U$��N��@Ū��F�9��ȎƧ������Ԕ���ˇ3z����F��lTU�X�aR^)o�39��Q+��c�q�顾��	FJ����䏆��� R��86bZ4�
 q��.$I��9N�#��KI	6c�ޒ�8�B�t��1��D�o�<� �8��"�EeMEW-���] �D1Ь��/��Z�6pnv�j��.�=ٟ
�B��@(hx�zt�E�����p�tP�߻��!ma5ѿB�6�P�h���Z���y"�w�v=�M1��? .�&6�yZO�L�0䷱�`����N�q�����V� ܴUb�Ŋ5��@r�E<�Aj���O7xy�B�!V�����=?c���N�\C.�����2?���ɾE#��L�6�%�=�<]7�ۢ"����e�o����\�3��Υ�8���M"�ߗr�z�u�{�r'ʶ?��/����;�	�.B�'ԣޜ�Yk|(�̲
�v�H�̥����q.<�xuŖa[_t �x�N�N(Sc�k�������~�Jq�PN������t�x�4�m�'ݒ������X���1Oe�\�"�e��O���
uϩд�vajU�λ��) �U�`����^�*��3�L�4:L�e����PȂu��"$>ȷN5S����$�@kFRp��)cah�=T{[�3b�t�m,��-����nA9i�/�|~v�n����-��z��&B�A`��/Y��\�J6(�ń'����a!��;��s#�E�z��Y�E6E4�]�c�?�I z���}��V�/]^�~V<@AL��9yS5��3���F�_W�3}����6�<x�����v�o�VhݒQ��M83�u�d��Gu*jV@�? w%��W{z	ici�t��Tf4ہO6i��<�f%Һ���W�*�pC��۝��D[\�V��W�3��H�C㻃��a$���	j&�.� q���9C^�7������1&�i�Q (��68L^N˚���9����oV�U�0�J8~������ΝR�!��"81�o��aa��V���2O�g\!�d�����a��b�O����ouXӖ����E<F��%$�Y�h�O��(��*�ͣ��= ��.���@�]1��WS��쳝z$��������Ϳ���|1QX4\���=�;A͙/��9P�U��l�9�x~k/5AN8���A��&�K2��`i�j�m���J�8�U$�=8o��������>Y��ï6\����C̈'�-!�W�x|z��Z�8�uT�w���>p���;��t�b��Ge��^��JY¬J��&��<��B��S���5Q���jJ�x׌�bJrP-hE�ý���;�[:���
��#s��t4�"��RU���A�=i��v.^�+�F�x������_���
K*��"��A�2k���K��f7��E�La���8r`>�`����m�`�/D���	����XȔ&�Q���,�+�(`â��Ng�+x�O����+��XO�VY��9���?��w(ڈ-���L`��x�lL���y�%��ʠW���m�$I���[��7��j'b��|6�X~�̴H��̔x��)1(�	��-��	�`�<������Z4����uǺ�e�7}�\�i�Y��M�F�P��]�^֥[��G�Wv3U��<F��l���>K�h��B�˱t�yZ}��n�)���ܶ~Z��0nB��-�Cj�^��Zb�-+�AE�w ���E03#5C!���%�q���z\71\�a�����0�NI0?��ɰ��Lw/�3Y��"�BV���E)���#���WQO��Kb&D�Y���(<�=:h�@gX�^���}���Z_
@�
�3+��aT����l�4ϒ�������_��sE% �yTf���)��T��y/8�%t.�hRDR�Ϝ�s.U��>���h7O�̜���A�)�ʵnXٹ��K:��ǷlD��v�9��6��3�	Ԥ��[���D���Q�i�G��z��`�	�D;�u�S�!��8s[��6ۻ] T�=�r_��f�E,�a����9�u��&�A��\|����bǉW��b,J(���i5b(�;'G�0�n���7A�Nt����PU � �U�F�s����/�y�4�;e����'��>�t�aEw��6Ⱥ��yy�K0v%�?�C[y��'��)V<�[rS�`��%ä��{�~�)s�I{X�'�2jZ�35�%�>� "u%0m_�����Q-��?$�kO�y�)������6|�]/��4g.�E=!J�E��0k]?$���ʊ�BS1G:�+�ں����v:�PC� >��r�<�߇\>3���ʉ���`'mmb� ��z)�mF�ڌ�qL�m��w�T��	$|�Y�_M��G��C�ItL��yJ5F��*ŲY ���{G�$h�?�'��~M��)3z��~>�hjR�?Dˍ�YhB~�(�Τ�y�%���]#��6d庣�#㬡���yݨ��s����E�Y����2/��1�э�߅�-ˈ�z�g*O�}�x�����q��%u"���%�B�j�1��@�h�.Q�%٪J����{`o� ��g6�:��A�BՍ��T!���/�oIq2�~NXZo��~��	��"�:�zi�7˨�,Y4|*���F�1����e���CŹƍ�ZH�#��:��l��y��*J1�n�c)�\~k��roKcČ�T���������(�C����	��n���C蟺jVӹ��3��>C�EFqWa���n�y�`�����7Y�')5��/�C1/dt�nP�rHn�3E08C��A����XY<fv-�1���/��t1ʄ����~*Ag
���bt\�ž+��n���G�`)�QV?)Uxn�B+u,QRSD��N���D��q{aS�ٺ�%�4^!�y\O�꣦,J��&�M=����'u�\���isa�e_���/�C�;g�P���FPϤ��4��� ���z�q��!�۳�y����%��4\k1��0X#VC�Lv�Q�X�e�'� �,H8}<��I�3�l8�y&/�>L�x�r�f���)1���c��ŏq�F/�A�Hc =͋W�����'��#����7F��BܻKgL�_��v>�X�^f��s�����1�� �V���v������l|�ȦP%��Y�Kg1�١]a
�7=,	�yF	����3Z`�G7�J��t�ae*����Y�.���7��m�����	T���Z�ؗ���Y�]z����A؃^��l*�n�?>t�Pȣ��jU_ ��Q����&��<�Ц ��$�7�
��B��������P0�@~�����M�E:�?6�<x�h^�
u�6k�ୄ�2(N�̀��������ΛI#��98���]/&Ԓ�tp�fֽ��dƯha6L���(���Zr���WD�2���O�^�i��#�m�$��;,�Δ"��NѤ ��B��Hd�ʈ���)��,�ͦk��0ι�q,`��p�q�.okf�a]/�|���,ۍ�u:�s���4#����?�*U�E� ���0�4�L¢��VV�i2�rl�]���E]���0�[d[{i|��';4�Fh�s��׮+�iQ,߼���_ܷA�Ξ0��a��
?axu2;xRcP���ׂf��#�$$�h���+���s���nCG��h���V�}7����<ġ�z�W�Nw�{� ��{�|Y�=79od��ÍV�=�\�f��y��Ƨ�|*�L��,I��CB�o�������`�(�U�1�@�ٹ5�y�GA{!+3od}�U����X����-e*w���$�V՘���Zv	����^ܐ#��	�6��:"�����-�,�E1Vћ�#ٍ_�6��lq��\�p��f��z��L2l��x�L�w��*<=�q��]����ZBG����U�N�9�� �&�
(Rt] ��s���|����^tWk~���/��I�/���?�N�tZ���̭O��;Z�'}���yP~u7`m�ٶ^�!9.�Y{���<�2�0#�S+w�%��p��FKYq�E׍��U���>�����Xw�V�JQtű������̙B����I��F���~��]R�=���+�������$a.��� 8U`���2$���ޠ��0��!<�:/��skk����F
��7n���/�U�4�=|��v��8R!vb��(v�s�V�m��j�c�>o��VkIM��dd@�U�RV�- �b��	�Q9��/#ӊ�#�R���}ѕ�zM򘨌��h�������-���V?�������%@�z� ��<�r�t���|��d��B�j;�]aFaI������|�?�ڻ�����
��4~�/q�ڵb����������;En5ƺ|Io�9�R�Aab�H�nu���xU_��b�.�N~�wн�+T�:��&o�At�2� �@��@�\%^���u�O�h1�ܬ��y8}-yW�CvD��*FRXdԁ�n��I�-Vc����w�{�wP�`J�o��'��b^��XǨ:t%)����B'��<M����6��j'��잡(fs�P����s��q�ƨv��$H�����Iq���>{��72�{j���CU�M,��Y��v�b~ X�.
��d���?�e3j0*ŧT87o�U<�e2�vO�1��!!5�E�����E>��������� n��f̦���|D��X\� �~�)[�!����f�d.ߨ\;��0��e`�:@��n?�HE�6��sZ6t#����7 �\{_��kH#��gS?�� ǜּ�Yķ�~��Ρ�
5v�9�1��[���BD��%��F�����R�22�3��$�n36���/�k��oO�D��$x�Q���* � �F�g�*zbM��95�K񴖑9�&�Q/�|Č�AXRoy�pY	C����L^���{���gUx��ʞj(E��o����r�^xp`G�ϊ☭7d���+n��/�a�i�:0�;�Z���� ����@h�,?����-�Ar+N$�g�N��4��)烼�SP������e��+R�F���ь�SȨ=�'l��$m
�@Ty9��#��>HTxч�`���~���Q\ދ*͏��g�d���="��[��/����7M�������E�'>�	�u��H�(?�Ao郪��[Q����#J-��U��Q?�<�=��լ��2�"#�Dud�4��Uv�tfvS�욜��QL���� ��B���
9��n^�o��&����]�n�s8g-¤�G��
����8Wq���К<�B��Z�U@�>���{���5�"�+�ǕR���Z���J���S�[~�@���[�>�=��&��5~ �iJ�VF�)�{��!�zY����5
�#�0�� ���k��?��Ir��n�tR�l^`���k�53>u��zv�yH��6�D�ܪ6'JmZS3|�T{^C>[L����%F5K+��Cx<"(gН'	��(��(�w�&I�7k*���6DD��^��DV�&HӬM\��s�cm[�"��u�,W,J�i#�%\w�A��F@(0��[@�;�����Lu��(���d_�� ��X�G�wsM��,��l����w~;��$���B$zZ٣�9Ⱝ 6^��g
ir����{��x�`��ٕ(K�<<"������:9�2���3�w|ҁ̣���hQ^�t��ꦫR������^�Y^���Qe�g�%+_wC�5�j%�{��3ʁVP�b�q�	��L�����}v�z�+�k�R�*���af��5��@��&�R�u1Pj��CW'S�Ӆm�_N5Nx���Zo�]����i�Ѩ}��]�ہ�U��pԫC�+�bM����8��R�¦��+��}� a�4\�!�q�$U{Iw�dF�Q�p��NWi}�!i��e$	.T�F{��ggр�ǹ�)U��0��Ϛ������b�6W�M ��5���t�Rs��1Ñ���0A��]���2����T�4D��śE�Ow�+���+�F�[���-�7h��6J���M�)��;�%���yb��I�"�/oT�T���4�E�d��w!��-(>�����G��_�ҿ�q5ʶ:�9ب��K0�F�ɹ���5>�,T�����v���X�h������;�3��&꾮C�y���O��������qvµ�t��A1` �n>�xx�B�V瞷�������|.�[��'![�}�I	��ħƯ�Kn�b;vy�(�8%Cy�{��^�Ӡ5�IW��I7a �]������c�2��E�q��)�8�u˩�h��zwK-��"�82�f��|�"*
�
#/�����  �$^�e���2Ev�q%h��xp~����Ii�Ul�J����@V�~]����<�*"�e|��ʜo'��f��D�������\ ���~3ļPl��'_�P;v�˼�+-Yzm��7�.�l�U�h� ��P���+���?(����1,�����yx���w@��dʑ��Yꘇ�5n�m���fp̭���;��KI����>��;2g�=e�1$߰0EˤJv<3��,�ː�*�orJ��:��$14s�ǒ\q~�Cך-�8V��HμN�4�L�Í7uJ��K��`�&T�,�Sv3L)�:X�����wEn#�^Ne&����G</�='f��m$ͥ���,��EJ���@��RA�YV��cr��~{B�c�^�js�S�'����}���������ߙ �/�E+��G���ᦅ��[n+@���o���r�� ��)/?�vHO�j�?Uja����&����C�QJ9���k�!��bj%p(��Z_�f+AzG������J��`H�\�+h�߯��5Uq����?(�|�f8G�"f�ޢx�b��(8���i�ݔ0�<�#��	pAŲ��I|?��6��.#�r�7�K���ɍ�~���d!�^_�JV3�g�Ɔ�0�CQ]6+��ow��ц�}�lb������)�y��v�뭴�0ĚFr�5k\�42L�TE����黴m��~DT#5�[��9�\ut���_Q��^��S��#�Ogza��f�xg5��Q��W�4<���(�=�_���8!�v�IrA$h�-�Y ?��/0�-#�¸��_���������X/K�5VKP�X1]�9� ���϶�>��%�����j�Z��xX�cc��M��NtWx��S�U3Q�^��Aw�.��["[^�l�@Yg��:�j#MM�g�u����`<�UX��u��\��ѡfڪJ7�ݲqb`�j��ٻ�H���.P�����йD�W|Z�E���ߕb�]Y���s�Y�X���1��u�3��ƍ,c��$$�cG���?���W���a�=.�����G���H�tc�����V���m�σxX�؛I�����]C�.�F2�l�h�VU���"���Si,#�������yO�%`z��TS��n�Nc��a�u&�ug
lY+��u\��$Qg�������+�49oIP�x���2��w�`4��_>��x�`�,T�iB��5����������$rXd>��&P!���OF{�6�(P@�����\�N.�v�o�i�\�7�o���eR�B��+T:�2 g�)r�,e�ޠᤸ�/=��ª���UG���R��v|�h�Ԋd��� n4�w�"�"n]�����(�4�O}i�]b-(x�z�7	�����\.��`l��w��W�TܽSu��9è*����+N�pR�!�4("�t��#%l�	��B������k��g_��U7Gb����[�W�F~[[��2���WT�XG�tr�X������G�鎋����H�tN��MC+7;�q�>7(�����ji�ծD�6��U�W����(8uU��%3򡎗���L���	�2"���������'Ilȝ�B��2��u�v�K;G���F���p���0��rN��M�v�'aTK>������Ѷ���{n��8a���;��sF�� �<���{�|Ѵ�L�ȩ�S��7��W�7����J��������h�� �5�{˔G�j��CQ�PS&�.����u��Uə�]V��`"������:M.�6��G�м��W�A)���Uh5�[8��V�I!�dK��z����4>Z�3U�臕^�t�3���[I���ډٓ_m������^5���M�j�����V�r� x��'�}v�����T1����,*=1��uυ�'�Mv&��|0���68cDR�@<#6���+�)�%���1EX&9�����*�X2�����:{_�Y�!˥�}�c�iCCx����؁]q��
?IL�Rښg#8��1s
L��!�)�vu�_���R�Ҵ�î��^	�Į�̓b(f㵨K@z��2���.�Qe�!>���Zꩉ_;��Lp1Bu'"0�C���g��^��#3ɿ'0�M1�G�����I�w��Z�����D ��r����^0j��O|�k�����7Ѥ���=�2�VLm��k~�D�9�5Ӵ�|E��K�%4?����'���:ː#i8������0���(�A��Z�dx%dS9�9����NP�F� �t��9Yȉ-惆Ē��C(v���;�N��$�]�mĮ�ch#xB�㱑6Rə-�أڨ��t�^��ϧ^;�w���� >���O[-5�n��f��2�u�סOt"�o;�(�I��͕,����ay[���!�N����}t���a�f'��o���;���\L`�y\.�u<�CR���yYs�qr۩�sϷ�5�f�	��簽���F�x9n�]�?WD�*Q�W[��Tl2H�-�#-\��O����7\Z��[��X����KV��?��)�G*<k�j�ɷޒT
[f-��uM�+G�J�5\��{HHl+��" �������+B8�BKSs����ZWAˊ�EJ�\x-�����P��,��;��1t �M;܊��$yo��2���z���(��v����\-�B�*��k[�K�e��ł�$[R��ja ���~��`1�� �p��\#������r��rG{��y@fiHF��W�h@z�y�WY�Jf<R���EF�W��*F��=b��y~7�_����!���TD���o�S��E�l�!�s�1��[mDh�K�A�VcT��MJ�M�BF�B���?���;垂�ik�������8���.I
/�o紐PnI�q�`!p�t�G�4��h��%?pTe?T��l�7ݶ%k�z�f!�5+.�b���ͥ�zb3i���C�33�zK��4��wx���Z*l���A��s��o�QS�H(�����MvH<+�&G#`�A��x7�ب�@}��0�b���Al2!T\H��U�Hl�2՜=N�O�����D�ϋ��׈�1j�� �N-�P���n$U�)��}e�ݵ<v�_���#uǊ!��@a�:��7w?L��}2~�/��q�fSk���~����g�52z�l�{��; �����p��G�\6+瞰jO1�Y�c����)�$��t�H�R��^Ge�T���� 8%����-�n&t��R:�zV��5ҁEw��îf�>Q�✢m���l ,�=�����Fn��������[0�_6�u#;��ZL��u(�hVA��|W]&'��`/v.�i�$��1�
�Z��d�?�ͨ���'�P�unc %|������R���,���F̋?@�R��'y���(��B�G���rmJ�DС�ݥEC�/�h�u�	��!�]�)����$�aM�B�T�bW�4Ē��;r�g!9AaN��|�4	��_�&P�o7jpͧ`nh���٠~����y��tw�D��Z��ZkV�rD/��$c�w��� �u�i*UR��8��E�OsZ�y@�ȴ	9�Q��Oo&����Ak��]li{4J,�OK��O#�"���3�+�^
d���X@�tg����PnUm����MoE�y��oȕ��G��,(����5l�)t3�vظvu`0��ߖ�	�n�z�D�����-Ƅ.$M��y��L��
���{S�I�����@{3��0��;_I
,�/`Z�u�nbS`��v���F����wg�K��Y����T�gVW��s<���4�t$?B:���g *���D�Q�ߦU�*fA���t������v�2�#k+��L�N)�B�-SC�p+-5׶?C%F�ܡ���i����@�.�� ����r�h�˲���I���p�2C|ơN9l�e�ݰow�a�}�)fű��q��.*�OLV���4:Ҏ�+h{3P=�M����(eT��'����Y'����Tx�s*и�q��V�P&�8-/��Z3j��Z}I�����������,فvf���}�q#1'3U����GN�>�>z����~+,z�X�n��"ħ��rB��%o�l)�jVwb{cTU�f�#vX'k6�ziwu�$���n��;^K�,��zu��%�٣?}�` �fp��T������}�����0�]9����s�>�AŘ�t/����zi��{I���Wԍ&�t������϶wwwl��oa�u��ցd틌t#��o�����..J!?��+�]�by&��ҥV�K>��0���Piר�� �Z!Fc�3Wq(�=?od�a��H��Y �[دj���K6�`ڣ���"�}N5T�ux�^'4���wEhE糣�YÁ�pڻ ɛTS�V`����=�z7r�Y؊j��ɥ��'*&�oc�L�eN�@��!�?I�ȱt�3	���X���mIX9�n��뿓&6c���� ��oN�U�ì�K3�a���3��0��3�Ki5�81<|�D{�sTQ(lu�K���n��`�BĘ����vy�uD�ua}S$h�-Jԟ�C��%�D�/-��R����9��z���311�i���T�k�Ĩ��̋��s}��Ƹ> �����ge��@�2w�����r�%2U�|Zo
�H$`Re��K�~*RRl��g�Z�Q 1�&dn��Rg6l��|�n؏����j�y}f���њ���!��C��Kax�Խ��I��J�S? �HҥOB�=��gQ��N�
25��_�u2��1�ϻ�Q��2��AH�TD$[v��L�(�}�OEM����}QH�f��:xO���8��;:e".'{��ʀ�q�����������f||��0�I�.Q_z�9
�)�o!����$�M�썩{Ҙn(i�V��k����(�q���{�H��1�t�5CT�����k�l:"*?��u=9�t�@�$�3���D������ �/�I?��FXC����qKR��_�U���T��i����K���\���(�s�@�Dl�:��*/��"�'w�9���S�˕��[f?�aJ�B�]=��� ��ye�!�wwֆkU���rn vjഗ� /Ϡ�5N��	Md˿a7���Y��[�x&�1�Q"��y��#w�>LsCbX��/�*7;q��qx�=Q�.,����<x$�`�?�؂kߠ�.���7�KL�����n�������㳗�����f���*)٢x�t�
�|z��h�m��K&�U��9�6Ι�7����Y^v��c�{�M"E%E฼�T� ®Z�����<UG�C�=o�4�)��BһlOc������cҺ�薚y�1um=�4���$(U�����;i�G �_�qMJ*�zq"^%�l���p#�NÏ��F�ϴ��n��zr��1h�Z�x!Ɩ��i�=#���md�-��'B��ii�+�T���:q�s��鳗�^״K��뷷?%�9�ϖk�l ՘A����F n*5�L�A�����$ae.����f���e�wȠR@L�>z���Ш��0�M,˺>�ƿM����j9�����-`�nx���.�v E�ː(��^P��enG,������թ�4�oh�A�r� �	����Y��*�(s	Lf�r{]���S])��zi�����V9.N�bW��w	gL�vY���k�0����w�[�>�� � ���Rg�⶚�4F'�,��r�3�)u=@ț��Յ�E�HK��0�Q�*�g����Ni�Z^}M_2�L��fJ���Nކ�ib:�@����%	���"���4��r3=�����'��N����e��I�D)�`a*�V�޷-���e�q۟�me�
�{x;c̺+��j{�m����e�����>�R��j2�(�]YJ⚇;J�X������2�yG]gŸ~�vj�c(C�DcX��`���YL�؂n��#�Z'KNV:o�&�;Z��!�f��H��!�����@�S�rs���qux$� s��
 7Pҥ��'�v�����y�+�qٌ=V/e'�,3K��8�������|˚�����0N��	�ܡ.���m@�mH�1��TT���n��h�����⇼�_U�e���Z��h�u�lzs��|���tA	���z{�qH���������W&�.-a��B����j�	�9d!°�+�z��'��*|5d3�R�2ҿtK�~�?��{��՞�
�M��3��\���ȹrL��,��y��R$���<��(P�4�#"�i�;s������rV���Q:�%g=A�<���X4�1c����Nl4)0_�A����9�Z��9'���mU�Ica�u[訪��0��d�\F��l*��Zl���l8�?+��8d�s\Q<"=_���`hClx�U�/���1�}�9�yDxs8Z�L����r���ooU8� �EIr갶�	0�tySی;�S����?�Go�j�;[f�3�Ё�g˪�nSe$`@��H��� {��G{����-:��=iU���V���m{tY���lI&�'�5�N��z�z�9<��z�V�VU�p�O�g�T:�����ݺ��VGϹ��YDO�2���O�����6�k!�W�in7�)[|T���E�g��gU�u�4��˓���:�q���?�{���{�ˡ)��#��KR��e�X���ݥ���ŧU�t6Sm�p�!9���,p�ozJ\�8_�B�?���(�{m��&3�	T�e`�rK�r F������p�y�qJ�W7�g���5G^����&�4AϷ?u;WX��jg�$�ʵ�j�M�]�s��XV�8?;�y�8Q��l���M�������`����ᔁ����,f�z�/H�����RPq>w��oyV���b�Hݥ��t��"�-�w5-�����ZZ�,uڮ$��{��jq;PQ~��u��c8��=�~��	�qY�ٹJ�>�VLQ�)����cwR�i�32�'_uo���Mԝ�P7,t���甾��un�L�-���Ec�`��3^]�e�:o��d�N��I�2ND�0d����L4E�����b�`�f�����;�8��#:����
c;�Ni8K^{m>�U'i����P��cf꩑�0ހ�/
n0����s%�,)r�%L۾�kѮѪ,w�=����=�)}Օ��1�l<GB)��O[���Rgcȱ��o�
�B8��f�`���ķxg
B�`hu�`M�h�����bH/T���Q�q�����l�x���X����Ք�7KE���Za)UBzO�~�K�#��)4
���ivT�U���#����D�!���
.(�+_^A�k�]H@��ݴނ��
�qS����� �$J�VV�Y!>�Y[�R;��y�L��v$�v	ٻ����jI=Y�r%�����h5�r��gL�>��T��U�_9S>��,5JV�����[���Tm$��8��K;����K�/��( d��JG
]z�|�K�,W�A
A|Vŗ�h#�U�z#UB�H��#�������D;�&��Ur�1K���HJ�]�&�0u7㼤�e=O�(	ȑ(g�ܬ#ݾZ��xG���������O]�^�l�ܱ�ʧɛ��1r��9��N���0 ����e�븮�H1���l2��*���6���x �ݼyJj�y�W��4����ҘPu8/G���0��� *��m�
��(6C���3nmVz����fL$<X���˜���d9�aNط�
2��Z`lN��4]�GQR����Z�cT/��,��6�l2�:�!\��xO�$L��8.�uX�7?�L:JP�Y�ُ.�c�~��A����r���+#q��C��jSzK��p���h*uF�Z�i9��I���8a'���C8�"�d�뻋�у{}�Mj�u����JY��� ��׋T�V��s�u�B`G�w���D;�ACb��pj�v13jos<�K�:Y� ��w�+5�t��Hg�q��*^ih���f�����h�.�귞�U��G����-	t�u{$[e���R@�:&��s%���]z����ZM�؈2?���u�?�7��S��57%��m�wSB�οD�Ъ��tg�K�g���8�-�ӜRw��b����i������E\���aaEnZm��	Ԏ:22H�>w�쀵��orץ/��_9�6�t�q�Y��:0��rU줢�jD������88!�ec��)�O�,�!(��`��Պt���K�C��,��b��:؊�*����6����x4���ٗ��z_�@C[W����؊w)�d��V��v;\=�1%.L^��4��2I Nt��RY��eq���`�	����$��0j�þ����뮿"k�u�}[
�^"F�	�w�ш��)��	-�$+�o�"� �B���#���%�{%b�֒�ѭߞ�k�K}�m���s����$`x.@��{N����0�	qjȩ:{�./�>�_�+�� �"V:T��h��ȧb��:��,␁)�^X�w�=��!?�j+ !�n^��9~��#2��$����p_��L���ed�3�u%���wZq��95��Կ���Ab9���I��IVZdčy�*u��	����=Ms6ʏ-2�<��۟;h��w�1;�*��Ucd� ��K�"��Ud���)��]u�ՆS����%F��f���/� �FB����T8�z��1[�P]������|FQ�V�����!h�����,�w�>�U���T�2����2��v���Դ�j�Ó�J�����x�u����iIC�H'2���K_|��y$˚
QJ���\!�A�3�5J��By��c��8W�J�N�6j XC�K��%%���k#&}��O�x4�Vq��-H����s7
\Į�]��z��Q�BH;D z�!g�͈v�ł��|���l����x�����ZOB~Y�9��)�C����L����g%�.�9~o�z)v�P60 �w[-ۛ-�����<��j�aJ��+���������Vb��`�C���J����!N�Q�����S�w�H�b�
[PsEE8����#�i|*�|���Z���7+�j�#j�Q#Pv|�ٔ�o��7��~&dN'����
�l��g����ȹ����Խ��̣�0T/)|c��
�嶖/�@k@�S��bc���W�X�6���0���?p�*d��]�$��W����'����ok�)×u�6���k*JU�<��'kĹu��Y��V�@{nɵב�,�t��=�����k�A�+T�D�$U�V&���B7�����=�괡��kc�8��5�5qncѮ������T�������3K�;����Ձ�A��N6��Nn%�����ƌ$��:�.e�}e�s��L��?i��'�<l�r;�o�N�b>"��=�`R�d���0�~�>މ��o������ĭR�����Z�����<B!RS�J@��M���q��ֽEv�݊�7T������
�T�gS�':���1�h��D�#�ӑ����v�c�}y�Ҕ�K/g�����$H��8�!�4ɪn��gw�&������bm(Y����W����T]%��[��\�(e���t�c�k��uP�``��o�G9�H���; ��*y�]c%��R�s ��Y\ώn�Tn���<p;F" ֝�Y?���zs���b�0��(/��D�Mճ��^`{U��lW�\d�1ƣ�B\��+q�&M�<������#�ڊ'<��f�ky�h�HN)�I��m�(�>��]	T&�~�5��-����ʘ����S)���M��r}�Q�o q?�ٷ{�����X�t��U�]f�Xoyep�k��<�����caly�1�ULg
�G
B�	�F�Y�V)���M�GAh�3�e����o�ZCx�MC��L�6��r!#7!�� ��A�v��QS�����	VJ3����><�.�/�1��I���<��	��|���%���\�d����X��v�~7Z�?|g����~T/<�[����fzI�Ahɇɛ�T�C�����5?}����XՇ��2���)p��'�CeN��%}_���'.�Z<y�*a�B�	7����ub^�`ɣ�̐=�d�%_Nb���;*���7��u�Pj�1�`��ֳg}�s.��CT�p�l6@���{�Jj�D��ȳ�!>�@Q�N����9�	"X��h��6���E���o�����pRqiQ��j�2�&r�C`�)��(�+iR�i�c�[TJZ�k�	���i���Mі@M�ɫ.=]��*S$����g�ܢ�G�a�x�Bn	���2���*���(�������1�3�C�����Tō9�e|����+�H��W�#�>C�p�F�������V0nf#��l�*|:?Kc�̂ ��g��(����r=�x��ߚ�<r���v��ìqֿ��/��8ᩆ��(%���'�Yz��`ൡ4�'��DtU��a�X������W�,{a�u�Rr�+�7 �p��˯'�=��]��VC�<��6�׎���$Ÿ�&�Y�Za���=�]��~Yt&4����.�0e+����ҨU�g�5�����ei��w���L�Aze@I𞧄�����'���x���]B�{7�{�N��{ �>�1w�r+�v`s��c{o\��,;{	8�#i����fV&�!YG����T�,����y��p{�ѷ��N~�I�9�p׀���)9�HzM��E"��2w� 1��bG��҆�k#dCˌ��?��
�E(q�]�l�Fꡲ���J�+���>�71~.�[eUm�'
jvϾ�r�I�#F����l�H��q�Qrf{Q�ǉI����+"Ћ/(��ĵ�`چ;,�	2ɰ���3��s�ֶr�.x���Y�Z�C���7�⣚����A�2�a�I�����_M<���b(r�^	��<�@&���kQ��IO<Ccnfb�����N���zdlK��Ni;KrbC�L����8`&["/}㤈���n�n�U�3�o`�k�?���.��inX�A,z�8sw�q�`�b8� �!��5����P���(��� �u�7ԘT���_�$y�����Y��x㮇�QP
�p䂀��^��<9C���ߤL���C-�CNc#f0M��m�"U�,f �LQ��AW�\?�#Y���Tqֺh`�D���u'X�r�t�ԩR�n���I���!���.1̂VS������*ަ^�N�%E�C<F�aU{Î�kD�jQ%����	J@e�!�ˣ�r����da{FK�y|X��M���g� ���%�ιqfHS1��A_o��fiq���A�N��D��fŖg�P.��1j�O����ϴ��\'���9��&���C�X����P�-��Ĕ�}m.u����v־�<�f
<J0J��t��f$ҟ-�Y�	��:$cϥ���ۤ�,��㤂�jO�g$`S������+�
q��⁎�b!D=<��e����(���~j��w����qE5lQ{�UV~�}b�ʠ����'\��?%�?��O���Y�1U���=�dZ�V����y㞚g�?q��4�=��c!n� �[����9��UV�vO	0Xl�8��[�� gWP��%�zM����e؍s!r��+m����QC�4W�1;�c��m���v���hړ�u�ɐ��CC8�>��@�j�L�ys\�_+�Ӈ�B�J�p�)��4�>����e@��B>�����$Q8t���1�Ԋuh>!��@�K�>>�G5��|3���g���-�#��f{����زYQ���|Z��y��J���Y�0%�k#q���5��'��@rO1@*}��6&_[� g�CA�V&4h=P����MJ�~��q�]B�S7'�<�[��6P��(����R�1�n G�v�k|��W_��N��^&F ���LL�dę�F�`��"sL�����E2L2��2���)c�<+�p�1a�8�*aak�K�4�#~�O�Zh��H���:�/�hr����6�?��џ��|��<����	�@{ą7~6��+E����ǋ@���R�~��h���X�UO�M�������d.R�lV�h��Z�4���z~ܔ��4�ٻZ �ĻF@9 J�B��@D��j�=�9���A�Mo�ݢu�=��A�US=�����2Ag��I��_k�}+T��۞�9����r^|����&1�&�}ް�B;������d�-��(2��*�h�O�<o����.�g������i��AP��!�e)�b%��	q��0�)R��{��	~�~��y�=И����X��V!�o�Zr�ۯ��L���|�i�)�p�{L�F:{����O0_Ғ��抠z���9����6����I�p5����6��>Ro,Ɩ�3�7��Z}0Ъ������4����Q�>X����k��s�f\��:b�u��t�Rv	S�h��O��n�%=遹ZWw�H7��8,LǶ�ڄ�����@3@�Yv.���V�py�H	ؤ���[�Wa���'�0X���2��@2c�[QN^�E�k��|�$�=pٹC�7�`w�FX�V{u̝ܙ���0OVv��iƭ���;'y��k->����sܬ,2}��� DF	9��T�b����X���g���Fİ	��������s���D��:�y�u9E�� |^Y����sV-#���ԩ�����KSi��.�
�`���N������;��ڤ|r	����X��Ꮣa��h��d�<k��3V%$P�*�-��~��W�/49����0�H }�r���/�%��m��d6$��`q'��О�8���ֆ��i�F.�_�,�)h����K�ơowz��K�P�T���R�L���鼯���� ����	�o�_$a���([��9/��H9�<�[@�6��F���L���Y�#%���0i6MW�"O�%�h�L�MCcz,aZ�_~�Ľ����s�e̴݅ �샛5پ���R-o��m�Ej(u�"5 S�2򦱮S�#��)\��F������-߁�$���;rL8��RI���Vt���{^ThQ�0��!�?��so���Nъ������K��R$_9,i +1�D�>,�J3D��s��h�_�V��j�窚����I�$�ս�f��� hyX|`Pkl�eN�����}��j��Q�j��[�]_�,q�N���?܀J��Ft+���jԳ�X뒒ϑoC���<IE*�\l��u���z\�#�`�3�|�*� ����n��,�@x}�$��=�O��(�!�Ι�>�\-�[3>;@s���#? ��w? x��b�D��&�N-"��i��Y*��ˁx�;����
(
���8_0
�aҊ�O�tJ��_�dn��M�}l�+����T0:�ފ����Y�ݭ{����P�]�TmIW 9�ށĲ�@sǶ�Ӈ�J/�yߓ�~�@Q����ϥf/�IW��1�׹4�1@Nm�Bl)�	f3RZk����(-8E߀�p�)�gc���g�SeX4K�����R3������СKW�${�{\�@�u�\��hR�Бˎ|6g�j�%W�J�U�N8o%9 ���m��h���?�cd<;A��Kߍr�J�
Q\E��|w��v	�����w��Cu�#�����-���3���Vk�Lg�fDS��O,:���?��N9�5u!7,��@$n��b���$�����:OҶ;������%Q�����M6,q�"��;5���Î�~�������%O��lӧM֊&b߅C����p�N��bA�;T?��c����`�"6����бm��P�N���u4�<8C��ڮs�Ri`�b��ɵ�G4��p����]���@�1�bIK��h.څs��{�+�^��ZT�)mW���''(�!ŏ띳����	�l/i>R�#�}I�P��7mn��xG{^��5�~�������Y���T�8�*����s C��R���UO�dh�Ԑ[��L��`���HJ&�'��1�H�Z����6DIϜX�/n�wF[�����?�L�Cp=��L�i*Jd��Ho+�L6�݇�\㧌X�BW��{�^��?�L��j	0�K�M�$G�<Fb��xzN:�|$��r`͆`�vn#`m���Ԏ��d�����������&8~��kA��F�z;��nJ:mէX�ݬ���^�.\�4�çx�緈�l�H�׉>;vZ���WR}�T�a�%��O�׾��_r���+��"��A=ĵ N+����Z��QU�k3b|�M�蜊���َ�G0&m�nN��ϻi�	�;sf�NSG�՗�lK�|7�x�y>�z�ɾllsU�1N@{���˥��T �+pnoq|q"�������(|��o��({����b^��F�ز��HZ�lb'���_����3�}���Da|�MAs}��y�/��V?ǌpi5��>�����=z�{���ǒx:��J^���@B�&.ޭ?�>dd�IX^�k�r����}��}} ����?�
u���{�a�o�n�?VHA���+F*P�-Ϡ���ٻ�z�݌*88��'�&	�Q�n`|A��K���#Ԭ7q�u��EOuLO�͕6ϯц�L/I���E=ȋJ�f�	0��sc�ߋ�N؈��æ5=��N���jc�G;"",J��l�V�G�~q�A�O��L(:C+)p�)nYHt�010
-M�OL�����s\��Ao����oFzK�[��rSS2�La!�g����Вn���xHH���ܑ�Ǩ�	��'h���%z��.�3�g�}B%7�����U�w�I�-y��T�kLM1���aY�~0�҉"�f �;~�4��C�#d��C�h[��]����2y3΅�=�l\m�&�3�}���KP��������A"�����������t����%N��Q����7B�2LLt�d<���>I7�_��^MR��2�n��)[�~���*ΰ�T���O	8��B^��3�,,� ����I�,fﰎ���j�S���8��%�MTa.f�b����d�s�Z���G|1O�	2r�Tl:;��W�A!�����N	�Y�^�<t�`�2(~v�差KA�~^R�mY,͂w���Jů%���ݼ�֯�	�}x�')v���A��(���1j��/}�&���?��%Ҍ��>}�F���!%>��ir�X=s�6q�-@.�g�a�`}d�r�6Y؂��|�������{D�tV�F�
�%�6'�Z�~�y���T��<�`ע�]�ct�]�*:-R����hc^´�@��Q��ڜ.Qi�����e����%f�Ǩu��Rf���������gc���_��)zk	��F��)�p�IeRe�����XR�D��r�j\r�*�/(e%���j6��}����X���(�V!�@�6Z�rT� 0�������~�DUXvK���̑RDa�>�e�W����FZ�q�s�G��i	k��XO��B��𮪁��N�w�;���a�âi���B��z��`�&�L�t&����h�f�2S��i�Ѥ�Y}C')Y�:Y�J�� a��PdW����<��|XLKͻ�2'����VK�`��V�f,'�pϼ��]�Mh��;���I�䒇`B_�i��8~]SO����1Gdh��)�=�	�w��qTg�2陱�Mq╒�*��� ��b=a�M��y�XB�$�ۀ-���A��`F�dQ=�}��J��k��)�y�FJ~�=��̥ld������we���\ME`$%=Na$
���,��������r F�d�<)9\��c�5�s���p���D��L�à�-��0:v�I�B�n?��c˄�E��Z���U�",�r�:R0��\M���d�6���/���GX�6I��7q�f%3��Y��5�:͡(��9S�{���D�R�年�s	2S���exz\��#!w�!q�+�Λ�3Z���3��r3 ��x�h�L�*X}�^g��+vHtt�u}.y�2�=�N��sF��ҿW�۽��
�/��÷p��˲�z�����R(k�|O�
TX�g�ҹ���Z[Q�i��-�}����޿�}o���"bS�*�W����T�F3Y)�#���*%�q�I�P��-��Zq�W���;��Q�X`��^��i�j`+���	�GYz�M���^��3�M�	\���V��Np_��-�Lk ŤX�ZϏ�dp� w��og��P��Iج�|V�A�]3����AF��1������:/i�"%�7�T`���h_[\	�"b'��/4�>���+���3�,&��2ex�p��|y��~xpE��}���`�v-8�T��G�cm\�Θвo��9���pȀ�R�^cnHKh]��j�X;�4'l̨�m��IG��Dn̮��s�T���9\QӾ��rA��;2��@n+w��migH�����;3�)�B�`��?��v�S�:��Њ�Z>E�;!Hq�u��w�i
��.!4��,���<d#QbpX)�b?_V�G�s�8����!�&��'r��<��V�$.�fA���T���H���ϙ �~$��[�<��,��IK�I��.�56q��/3�&	��6<D��\YK�8n����d�����TH�e��lsf��t�L=����	.�� ކ�����J���L�+�y5�.xD��&�e�#n[Trl�Iܙ�^Í�}����ﱟ�ܢiƈ��iщw-�Rn�E}��ұ)V:@	�I7f��M��9��3\b�b�c������m�iޭwcV7'9�lvEV�j@.m���z�>��EV[L�TU��%k�}I���\ˣ��#Ƿ��Iҭ�7!\���h8�@�<���^Â$b}M.�|��u��ǂ�
0�5Ñ��y����[]��Ů@�o^){��B���v���n6��D��Dy��a��3n2TĐ[���P�Ϳ�eZV����8����}c��?�6���Y2"k� ����48E~���B50���P��O��-���
��uꛠI���?��d��=�3z
X|3�+�eJ���z$����O��-�/��s�2��d���,?�"/�fu1��?�y�� ��ru�b0��z��ͧO�6�PDv�Udz�!.v�F$�▫G��O�9��	�Wf�Is���Z^z/�wNsM 91��7�����8�gk���3Ww�1�h0��C!r��F+�T'�ɿ�j���N�4��E����h���w6��mz���p
P���X�Х`O�c��*s7���)��/�ۛ:�7ˇ�]aeHc1��j�W�!YW��w.2����h��|Qw��Q��fIu��ݞD���K�B�n<�ӑ?�m"��hi0��#7�~��b��SG��
���a*:�J�Tm���^#Ȓ����ϑ�|��d�ףf��[d��j[�\�`&�n��V��g�.�;�n�x�D���l3�gkA�c�P��p����f� �.�������-��)�3�*���:΢�.!�^��'Y���X��]u�D��Q�ΎE,�Z#�gw�"��L};<6ز��o�l���M�Z��2w�X8n�:�,��N�5��<��:��֋�~Z;��.$���p�+�y�J��eF]�dPB?�a
x0��X�*؅�pJ��	~4I����h���X"Vb�6w;�EA����)�تB�ri�D��3��>IdG��!�1�{w��; ����k�c�S����B�ч�اc������PD{�
C�:�%G�qV��A�&K!��j�/�=�os���V�.�S&�3�w�����K��(@���c����0����bldk����M����.�2��5\�{�l.|rw�E_�ݑ��7�zQ���V�?�*:���׋h�ʣ���C�h�a��Z�=��=���R�A��<��v�;}w��O(Ǟ�t4TPb[ow���ږ�pv���r��O�P:Z��u��4��2��%�|	����l���Z�&���<$�$�7�mL�ҁ�f��ظ
�I?7��t�Y��3$u%�`��� P�ݡ������(�9Bk�Ő�����m�\[�r�J��G����xby/��FX]M�OKn�p�]l.����"{0{B���s���&v�;���8PB�_(JR�W0����>�)��/�x+n�Ņm�D��2��/q]�eo]��i���=��
	R� �����		�~
":����f��n��`�Bw�0�hS�®��zF��(�(�� X�;C���Z�ւͪ����?"><B0��5Ǣ�%��j�;��D������ѧv�(>�5@�5�1~����s���uS3wۙ��"��bY ���?܎Ǔ�Oހ`����/����<��^:������[���I��/r�!Oۙ�z��
���*���N��?�H��Ӥz9�ҁX�#&�p�Yk�tZ�B�}�K��
y��?���ٵiSq�)��e�AV��M孏�h�)դ oCE[)��]�7��L�Z�=jF��O�M�:���6�@�Nfo0&�G��7?x���
#O����I5��_����B�u���p�W��E�!Ij���{/ ��`��
����੾�\V�9 ��u����;@�y94<�q�R�7ZJ�3�����ů���OE�Ч�^i�TI2��%���M�4WèU>���2~Q�R�%�+>�t���Tk�=���:�Ч0:K�pM`~E��[���׸h�
=�#\I��/¨���H
�b1
t\�������A�Smfo���O����m)|*X��N���p�t��kʭP�	c��;5>��]�kB�Zۺ �;ua��>RB��51�%����'tM�sH�t��Z�-��to�
����7�א�_7�-���1�rV${�š2�&�j!K��i� �w$�%�{µ��A���,敘��x��=��\����j����8�k��mǃdt&�e��K������'%J]��7۠��]�f�ZZ����頋uҊ����G�8��}]��'�mj�Q�ǣ%dqgg�6��K��o�E��#r������VX8^��Aܴ�T����*�DUe`m�;Az��S075�	^|�-@��M&�=��
���{D��0�:l����˲�����|��]��Z$���x����;�=3��� Q�n֦b��C�*�&i�kd�y:aC��;FA�N]��W��]��@[�ܫ�;*s�0��<1�n&�
�a��ht-q�^��JI�����N���ۿ�Z���B��}a�Ǳ��/!�IB��v����J�����Ṩ���0s �|�N1�3&.� �Y��'��e~� ��A^;�7��%�}ua|̸�O�V�Pԅ�GH�ȶ:Y�H"V<�R�̢�S��+h�M��)�r�?S\컇��M3K�;0�ʤ�-���O����ڰ2�|���#ZR�S�v٦,֯}�Ԯ����+�{�m<B*�RQ�wM]��@��yX���V�d�P}H�-��W*�YmUx��WdI��w� ��o�����*�D�%����8��B��S���
��
"��lI졠��A�}`��"��ʟ�C�u5!?�G��@%� l�)�;&�BH~�)Xy\�\��V����n�K: ٝ�4SE�4q)8�jj���L{a�'��a]0D�<Ώ��\��Z�Hu���L��~�5cGi��+d���OR�5���(4]��lf5��b�z��ߢz��Ur� z��l$��1b���r��K%=?���IH��@k�J�ʹ>����^�0洚�D.��
ѯV1lj{�P�Vw�귺�yp}NXw�z����劭�`�Gn�ˏ�̈́��K%3k_K?Z/>���jj������q��j�4B�\a���$�E$�c�B{�;����Q����z��"*��O|��^�|�Y~��~�2fD@�Es�{�@C�����x�v�0>� �=R��J���Kw�z��,P3�<CE�$��_�5w�����n�ŷJY�x%�����81�n��<���������E����kj����CNﭲ���̎q6��>��X�	��ŷ��>eF
�5��)1���U_3|ݤ��B^MZ�Ur2�
MZ�GHWm���\�/��L\�0�Mފ���Q���0��@}=W�J����a��s����J�^Ǟa�S��"�^>����9&��`�6��.��H]����i� �k���P3�yy�К2��-��=W�1�����Z��2~��A���MJ�����(	�,v&�R�ʫ젖}B|F� ^�
q�P��QJ�`j{�,��	����\V����|�%Jɴ��1 �Ӛ|����#&{�h���Y?�ڀ'~	(�C��7�c���/���zqe�����W���~,��An��@g���j����l��7dz�?��Э�P��v�	�j���m5�m�c����^a߄q���.7k���N |7�Pa���a�S1 7\�X��>.�l�2��gX6,�,o����������Q3'f�����z�y�b>Y�3Z�d�;<9
�w%���-b�lN�3��jE^����3{�%g���)�%:0F���dѺ�K�����:dJ��C��Lv���A"��k�䠶@�{��r��r^<�;m҃D��J�~+6w�`NyyӇ�6X�Z�?��<��� /�?����U{Q�Z�\�(�c���4&N�|i���Wd�Xv�k�V�1�I��g"����)k?� h{��(Psp�6��~0`�H������Vދ0�7~���J唤�Ɠ��F�rI�C��~�ei!Gb��[uL�&�<�	��`\����]-�֤�wϟV��W$�l,��J�Ik�O�,R��uy�L�����U��P�sJt�(JY����>�k��'��{��A�c\�;(&Y٠���:�t֭��:�wUO��&a�굳7��zr��+�����,���W�5@�[��%v/%�̞�W���W�U�w�@��˂n�ˑ;o�>��A��Ǻ��s��lB�ˈ�o(,P95�($�BT���0g����]��&w��
p�[j	&Ҿͦw�Ȅ���pW�2.X�ʔ@U�u^�E5f�w�wǪl�X�ߥ���������5�=ȸ�E]Nk�VxyM�rƨ��1�E �*�.���h�9b6�!�Y��.Չ%��"����ԺoL��rѰ�]�ٖX!�m6<9�XT���~ᙦ����@�-a�(���bŖ;pM�Ɛ��[�ߡmM����&�Fr8��>��E2@��ݕ~Q�6{	{QB*�?��Z)s�H�%p�y5�x3��Xk�G��mK6 2��
��O��Ѐ޿	䏂��@���xe�j�_|2>����h�k��z�@�QAh�Z�0ɕ�J�����4sI��!\x�W�P�ΧL��.i��d��%��ш�������G�I�����Qq�A����~nTg��d��~�?7�Ѣ��aL#O��I�F.��L�(��	@�Tŋ=�E��>E�#�����U���<�,���<QS2����P3�/(�tP*_ �Ψb����J�z��8㿷�lz����3B�yk�,N�)� T��&��]
^������n)��~&*/��d�������3B��f��|�P�ґ+�u���H�@E��@D_�է�KR���h
�L(88+�s#Uf`R�DR�/*�Z�0tĲ��u�v�%�
P4(�+{��L�^=�S�iUA�};V��,@`�<������Ϗ�k4�1p��f��'�fBL_�p��'�h	��03�O-���Wl;ɿ[N-��訹u��d)���$���G�'��-���,�[�봍,����D!7��b� \G1C��1U��D�RvF��Z�$騅M�o'�4�^ѮTw��B�y��̳h�7�'���9�����l���S�0��0U^�-�iٍW�-��.��N\�ӧ ���RA���,+�!����s��O�����I}u'�����)m�|��7�nȨ_!�A���I1��t��M�Bti`�q8\ݤ�H�X��p���e�E�T��o1]OU��H�	'���aR�F���j�Z8[�ӭ�n,V�6��R�����\y��
���օ7R�OM=�ܬ$Q��:�NEA���)P��eiN�.ل[IF+�����v�)��W�V�mlf;D�d�ؖz�&u}|kb%#��R��d���C��(Q���yw��`�T1����w���� �(�B)X��/Bw�[��5I�/����Q�*(���P�GQ_~�E����=�Ey�s�ѽ�ఊ@�u`r/�Y0f%Q�C�愂���D��	ѳ���֊E��%g6Z�*]�?3C��t:��[�CѸ�cd�.T�P��I?	�F��9���]�N��u+�f/�;;�	-��R!�
B�bء��S)�Ѝ�ŗa{�����X`C�׶/�\���������<̪�$��M�{����E���g��8���o���rs4-Uk�	���6��R�b-����LS�o���l>�տ���D6_�w�������.Z�#m������

�%6�I�]7�Ѷ�>����̖	�h�#�jKT|ݪ���\D3��W����]��}��y6�g.��	��, �*hC�C��T��g!��R� ��^�2�o�xİ�/�Z'.U�ë�#�~X�$�t_sܽ�
K�J�5[��DY��V5�OJ���R��v��s���.>����n�t�'75ŴO2s�Mb��W��h�}-�O �F��iU1�29����a��:_���\��+|(8��r�B?����+�.H��56w4�h글7C=�
R�0`̿��<Ѣ�� �o�{$7���>o�drc�6u��Q�fqĦ�����^8��:7f]�oܣ���K���'ں�WD��z�1�n�=ɿ%�`*�@Y���g�Q��s�},��4Gd���&5�B��_6�/���~t��R��IR����fխY�[$
�:O��Ό��̴2���,:��P����a�&oR'�Xj��:u�$�9�'
��Nn#M��?���^�FM��gv?���>�.L���POL1fD����9C����
��m�W܂�1���H����S
�T�vڈl��t)�����M*';��(��%o�; iWK1=���УR"juc�5v�\2Ɍ.&�K�ZC�e0�����~b��N��LW�?��G^�!
	�v߭��^�	�|��ti)���R�c�-��r|�u���]�Q�F�l�хk����Vxܢ��ǃ\��?v9W��d���{
w��R�
�I�� զ��
�@^)��H/�4�7�i�É��-/�yC��;�ҬC'r]�i�x|g<o�1�������*�2�<Nz�7z�-sM�{,I���03�Pyrn�0z��j׀��)h@���A�]3Z���xD>9�A�K4H�6I��y+�hi���n�[8�T���w��K��F�o�i���ߩxC�oM�����L�	�X�{m��Z$��!%�u%�6�<��	
n>P�ZLG��[|?6fmp��y��bf��.Z~�v"����e�ۤC�����J.�� �(S��.���?�~R)M˽k`��Qy} !j����hm}�VVlB����� ��b��@,�+�8.��ҽ�����r�5S�N�W���.3m����x|��d�Q7���u/G��F�R#I�/��� ��{�NW�r���x�dWܥ���1!�'ζ1_vC}���f���*��[s5Z����h�ҹ�����mC{T�I�7���A7:Ɣ+UO@�����m �Mc'�%����;������F�D��a'�P$�iR��6�]9����bg-䳶N��(��������C�q�R6�G�TL�M̄�C��#�w��gT����G M��2E�:��J[)ƫߠw(��ř(���R�p2h�m��r��&�U
���-��n\�g��Vì~8�$`�:O(:�F%T"5���(_������u�6dx�K�)��\:�n z�i�B�3�R)�o)u�,�-}֩i��)���I��*�?;�tĪ��G�w���{�?�
u0*$oP��|�Ԧ/���ƥU����h��*%+� �U��*�u��T�u��qt�y��������X�g�v%@<f�%�A�2�F�e��)OE��Ħ���E�pHY��s���r����ԕ�BR<Pg�m �R\��y�q����5~�E�	E{��Q�nΔ�Q@9w�^6�c�����Mp�2MK\�֮!��!r��B�b=� �L��98#Tw����I�yrJNh�t�-�= ���8�]��s��E߽Sh���e���O����"�VP��b��������j�' ��_������]��d�؍����Z�Pc�Y�}�,��3O��_���N�C�����WG���^���᳨9z�[�X#	���F�VRJ$�u |<�S�)�'�ʌ�����m���W������ƐY��	B���l�F�r8M�ݲP�x��(�R�Y�\���a#��k�ݨe���¿��>�*��ӟ#�U_!�szwKAz�ܡ����H���?�0�����OQ�B.go�f�<]��+tXv�?�t�~���h8���l"�]����j�I�zl#״�3&��<Z�fTF�@|�\��|�@���.1����K-U%����;�����3C��m����x�N
'�3��*����e�-�?i��Lv��v=��e�5��k�J���w+Nh�(I����p�ˉE�f�I0	� �����?�����^�j�:E��6�V�V��8q��������в�ϔ���5��><��ȁ&NP��h؜�N�J9l?W�{1��Y�_�J�D�QKƤ���0��� ;�o#����O1�+��fA���"q�o#!��8���&��B���T�`�_D(�L��q�%��3
�p��d���L�y��B��J�D��-k(\2�J��K���� ���ʝ@��e�ї!�7��L�9i��V��k��,6q��`*�\Sc�D�S��y�;.�W��E��VDz�-�d���>�5�5'<��B )v$^�Z��x�55xi(����ɝ�@T}�Ņ�]p��ڍ�g�荏R|y�N���=��rk�;�82N��ye�8�6��/����`�蟅R�K��sw�s�o�h�5`���R��h0�S��i�;1CF7�U��m��i�g��D{�4�a-4=�Us�osI�z-	�?.���b�r��e��IC�Z<P�qN�v��ن�#, ��>3�K�!����𢸛P�����4��1��Έ�,2�.1���>�<!�I�Y֐{��g�\��0c3��~��!����Mz	`��p�F��s�����dh�0�[s>)��4�@��:1�\Q/L"׻����L5.I��T���4�<�'��WT��cSo�Ǽ�5���ɳF����*�Α�e�<��8��S�D�o��o�U���/���9��;�d"�M�}7���4c�.�Q�u)]���X����_V��I��_KR=�`e7m}/������ʄy��'ÛA`��?�1Ƚ���y�`aX",v/⭳�/�3��߄L�L��=�O�Xr�NC��0�H4�����X���q�P�
)�����=b��wҘ3X��u h&��L�(�J9����܁D���/#)ܳ�ͯ	�vDf�R��8�D3Kv*I�م�&o�e#@+�ݲ�ǟ���wl�h
���g͒,�X�b}�[����>0�q� �nf�;��� ���F��u�����*8�m��{/�P;���y~�ݺ�{�%x_�Y�l��U�R��'*��V*ޥ]��!���u�U*3�nR/K;��Ch;�)K(o��t���"E��$	Q7�#��Ɗ�"e���t�m�C�F�
tī���<�'7m]/��
WN�e~�ƒk�v�7}�V��jÏ$t��Y�PR��Vh&����ҙ�*ǉg@!x!zs��+3\dʽ=)�
CX(����7���L���,�v3�4�\FGu�.��Ҝ3�?,Ky�b̺\4&�<H��-G�v�������1������݆���(��Kۏ��ޑ<��L�\�����U�����-�����~�a�/�e曭�v��˞1�k�w��x�d;m�C0���L[��Q#;v����P�N�]c��J�ߒ��TO�ۛ�Qm�>;h��|��񁜅~}��!��`ߑ��'K�=L��H�Ί`�A4s<9}d*����gZ�V-�b�v��.�7
n�9"XCNj8��uٓ ܭ1$:n6#�xM�E��&��,�;����E糱���<
���6q��@ʶ��>\I ����Qe�oZ�\�e�� ��P���S��_AC<�E-��^�Z���I�Ȼ�q��]�]���|�����,����s�� �ݤQEqw�<��)����w�7^+&B�Ox�8֐%7q@�-�J�x�:�Gֵ�H�X��A����_c�#����t'�.d�D��`��	�VmU?a!FE�S���6O��aNl7��`i�I���3qb"'%�nb-~�;|�)�-���Pg?s--�+���ϗW���]�[�Z����s޼��uO߹�6e�V�Z�9�m��4J��?`.�H�w�y��f��t{[:Po�\x����bM]�g�cض�5���g�E���_�F,t�����h[�L��8�K�7�=���\/"<2bQ��j����6 t�f���9%��C�ɧ� co����a�]����.a�ӇDc擽��/4K�8<	O��X�ܝڑ��w�0�������ث�u�=���ٿ^xT�WIdUt���͖�,�onFN�l�b�c��z	܍70q";P�[�0I-ݏ-��!���\�E-�N�j��m�v��@�z�"5%���m^.눑�K���r�wS��㓈Q%��x�~lB�8�?� ��@6N�5�t����+�)'�	����ν���FBb�P�U'�Mݿ�9E�c�-,��s{h�����D����S���K�u`�g"�p�5(�~�3�pɬк�B`QIJ
=��\�8C�1�Dэ�[�NF��|z\���\� �Ӽ�,�������k�o���Շ��si�?S��k�:��U~h-3.�`�#��la��vfإ���7�E.rIA>&"`h��_����}��Pa=	�&�B�&u���p�O��V�K/���<fSy�"�ZD�]1HJ~rO,�uNq��z�4{c��g���O����|@�lCZ3�v�8�'��Kg����4�<�8k-�s����nT5wT�I�ۿ�Yc�ir�}�z����'��|R�_~	����h��i���*���pEn��&����6Ҡs����jU}Kz��ċ�I��l��z�~�T�{��:``��[���F�Q�gs�,�3��Q������#2��z,���'�/�ͥXeV�:��z�(�c���NC��;㛻��Bb��.�x�C4�Ϝ����wj3�5�_M�/����ҡ�����W�w��A��ʿ[����@
�G��s��p�Ml	���_��ĨB/"���m �ѽ�T�J����o�n�b �]���Q�U����W�~�^��=�.�Ph���{u���ﱓhEK�nڭ3���nu�%�H�	�I2-ƹi�4�_9��T�f]�A���#�><ô�^�7�K<�v=[i�WP���@��J���e@�
#�-<l?�Or���x]���]�,�ɋ�cOH�~'A�x\��Y��sb���
��d<��rO���-Κ<4�u��Y����s#w���^;:
��g�t�Lll�;�S`����YJ�N"3�ip]aa)��=j ��E�������{���]�f��v����-�J|b�Zu�����{�Y$e���jr�G)Z[�P��f�6��EC�1o���6!�h:bx^�� �Ad!y1x;R �x/�#�E�-�C�T.���fƃ�h0z�0?Tqt�	G�M�n��jK�����\�w_�U1��%�1S���v��G<���Cte�	�O/K��M�1�]��rHm����.��5�����pnF&��Ki��n��GJv�tQr�<��V^N�?j�v!zHN�(�EQa����v�8F(Q`HǞ��]&��0��Q���@��F�(�t(,�2������H���qU�Pn\�0�>q\4�w�ZsR�{�p�G�M�D�C&�ߊ��R���c:����x����F)��r��5y$��}.Y���_�k��G�x�C���=\Jd���{�T�U��?��$�/�Z'�'z��{u�'������gMwtP��i�y���� G�js��P�<谡Ű��B6��l
��8�
lwW���쨁����r1�/�PQe����Gb{*/4���z���F��j{P�
�1i���I�m��H��,�~�"��ނ�I=���؋��a�# ���G���|���l���f4T8���̈��K7tΗ$5�e����h��ta����t��ۼ&�)�zQK�;�O�ȉ{�e�h�#�t�wz�>^���\��{���i89��(;��8(�m�Bl���<�����l����wyV��{7���=�%x�]:ÍjB��EO���(�-����h/)���~�&���N�� ���U��4DL�k�?$�<?��Hz�`fѳ5Cp��g�L"Hg���l�ĔƏDTx���f�Y0�<���
���lp�PN�WQ�� -�G�u��X z�)щ󺖓����R^��nBV��H&4�+>%V�D8ڡ5N�y¿����䞤��d:�JNG�֌��-�J��׌��`%��I3I.�1����(�E�'�1���cR�w_z�G���Sb꠱[f@�b�2Zdg�z4
̖c�C3aVwO ޠؤ=�b�!$�n�,Wc�g �c�*peT^� +QIv���(�_&+�!�@���@����w�p���	T3� IL���޹�L\�����0��ڥ�f_����;�Aӆ�ol�m�c�j`��ŗ��a�
1�S�+^�b�(��������Z�X��߹�����c����Om�����n��iL�{����'��u��<����|����$s�r���Z^�dt#h�m6�Ѽ�@e�z�����U���|\��f׿���V�������=�l��S��n�8�F*�E�E���,�������!Ku&��T]��_�LS9�q��&��~-'CĂ���9�vdۉvE[�����:��\l�޷шl�4Ȫ"���e� ��>���h;�@��.}�i���� qX� Յ��`0�&%�����m�g8

��q��f`t�t��yD�&ax���S���Ј3�m����3��n��kf�x̫� [��!n��i��獜X�ւ�幓��`E�a$+�~��(V=j��l.̉�"��q�d8AȊ�-�8�S�F}�(W����x&���aO��D9L���oEW֌�y����b�6Hsq�����ZL	��iv�������rұ�/j�H=��BX�0v/��i��o �C��|	`�Ǫ1�"5A.N��ts}�k9�$*��Q��J�BK��}����u�M�ܤ�|b�?�R��[+I��x���j�'�ױ��#9	8������ug|8,i�$���	+�͕^��G�w}����-�-(�@	����%�-$�n�����ɯ^��F9}��W�,���do#��mC½�d�F/���;a�v��/��Ri�®[�Њ��&6oA|��Uf�EȖF�Y�j��{���,��p�Ь���sx��ݪ��ȳ��ީɗ'C�O�� ��&|�H����1��_�	^����rEN��~�Bȅ�%`��9�[k��
f��\eMl�Et�)H%l�<)�dyXi��ܐ`Dk�h��t�ߣ��>��#�(4A�7-�$I\�.�טp�!S0�]��9u?����m-���Аv��}˩a�d\���\6�F��z�T{ɞ����C��[�b(�`����}'Sy��C4����s�X!�2��	�� ��jF\a�v]k�g)�K����-�t| �-��F��#�|m�aʴy�!~:!f]W�>+h�Ȼ�ߪ>׵`�U'`,�]p1L��堤�P�%4;Oǌ������i<�cX�ktSx�E���xsN]gQ^�+�.��j-.fIwz�?>��,,~�<0���6޸ �x?.	-�&��s����`c���ɋ��aȵ�CLO��������:0��5xTլry�ŝEN9#�tY����Vwյ�;y��g:c�k��A
���P��7h!� Xr[�N�w���gU��`m�]'?��@0!�@���&�7ho��!�1���4�+~�Y(>.�We�}#֒�N~!���_��j~݌ϼ��Q�|C\U?�f��O����MVT(�dր[��
S�tg�\�NL�t��"W"��Ȧ��T���`֍nq��8��.ɝ� h
������ �3W�\g�%n�FV�������՚�P"I;fN�=���B�r6�YVɁ�t���RI /�c���$R�Η�x2u�i���(���zAQ'^����:�(��f*�f��9�n+]�a���,�����m*�߁|��' �6fLgn�a��p�T"S�x�,1�1�$$����� gW=NT�.|���ލF�&��r��YG��&�#�t��cͶMX�v�K �c�9�}��]i�w|�!�gaw���*)���Ū��5���鱌�������V* 8�z�Єl��2xj��\�7_,a^��v�^lt���w�$��[,Ä��z%N��sQr���9�{N��_��>�%I���?���S��%e�]�	�ܟ��F�}����'���($��� ^�x~-�S�J���o�=�2���t)�|�Qt;��"28ŏ`��C���ig�1����Jg���!ٝ�wio�.��ѹ-.y#����|��w���d�"�r6P�k��yTw!o�x�Z��v�Au���?��h$F�+���3&�J�Ү��Ej�1�a��;�r��3.B�`;����ʘb��W���Wk��0�y��v5"�F������?1K��#eu��A��|����hԸ�hhkBz�^���S���p�s͓B�E�5x��'dLf5sE�2���In#B�K.p�����C��`n�3�Z�[��q��	Lh���'�e����"�e�<J�3a��'�+���.�"���DpH��c����|�1�6���.�#�nVh�k<��7�a�<a|�gI���TSkR�NO%���z��B�����{�|�[�{BE��mXa���/ l :�f{��{zx\�d!q�a Zd:���0@wy��K8�g���@
��\T�Q̞^���{&ˉ�['R#��~$���c�z�v��F0-gYJ�:��s�Ia�td�~��@��[(ɔ!�yM��{���r'gP��V�H�$�#ca��>tB��}'o���n��y�ݱ~.���W�׳�m�<XٛB���hI/Ɍ;�V���p�@�����j�sα�(�]�OeL�A_��]ĺ��6P�b67�W��9�h��x89ee�Q��QE�)E+��P �O�#9!�ͬa�Y��D�E��ۀ���*AJ��Yŷ�<� �K�+	5��K�*z>�����m�bf�}Q4<�J�g�qJ&u�Gf��r�����zP!��%{��n�n��־0D�,��T,+%�A��L.��6��He�r�ֿIp�ѭ�{،T��=�A��Р��w���E>>��P;���'���ߗ��ff5j&�?��k�G�8�q�y0�[�lզ^�LW����C��'�=�7S�x�L�@gѥ�Z�-d���7t�'2�a�])H ���æf��\��el�ev�|$ev��S����xo�X�^������yosU:���\t'�w���#���}ƞ�#"���s.������6��@6���z;�J�!v~��A�R+�#-o"���m�ӗ�R�l%������۱�b���o�\_$;��VQգ>��av�t~��t�(�u\Ȱa�[�ձ_�|$�������
H%!"�I�5��Z�Z&��,k:Q\pg�
p����I���N7\�����4���q�Ế��W��Dh�?z����Ԕ�O4\3ض��~��G�������;��W��d���#�V:N[a8q�[.�������kC�m|A���݉Em�^�;3#�<�P��	S�<t�ո��;ܺ�IINL��mls���wd��W�v�D�f�k;I�E�E#�wѧ���{�2%u|�<�*�B�y��^f�ӊ&�j��ｼ�FMC�d?�q��5QEZV��-�O���촇�ͷ/�����Q�%��u3{�CS5�2���� ��P���&7�c�'���:��3V����Z�����(��7P�I�bq����W�Y����?��Nz�#�*ܘo8Qǆ\U �U��ܑ�r����F��X<#��c�c��p�r��܅��뺮���V�����]?)��S`����}yaV��0M3ݚI�J�� �tα�����E�M%P���y#)[|��*OAs��
�h���o���(�� ���燯3NS�Wo��Wf�7,��6��Pv1�4��!k��G=IT&w�Q!�����=�ӝF�Dy�ȊQ�W���4���Cs��ˤ���)�N���S�g��^k�O)���6�H�Y�(
䒗Ә�t�Es�ZbQ��Л��Z�����\�;�T?ڝ�%���T�t	��:��:Q9��ܥ��8�{m�	��>����f��Q$��S�𝼡Q6צE�Y�L�P����l��4btG$���W$�}��,�R@D�|�4�`�(J�n>6��P7�(q�{7�����,eq��_�(�`;�\����;��aV[���R��iq�n5sE&|V�l����&k�i�O�܈��}�h�	m|A�\of�k<�_��;�K��uy��S�;]?H �d��x6/_k�o�&�JX>ĸJ.�!�u�:�����sс��zS�b�?p�L2�R����ʍ���&�q�k��D�>cB��� 3�Ʊz.NbT<�g��҇Q<UqpjI"8���W�����Lm/=�z�|�b��L֤�Q$R��j���qlm�vn\�|�������	�q>#(�<}����l|��_?4��߄COщM�:O�?����]�ĺ4�!�W��P�ўRNn�m�)�f}/���T�_{�j7q�QiN�<yc܄f�OW9"kR����RvB�WƇ��f���(�9�^�ʄҬ��V�ã0�t	2�ލe�p�ֶO� ����`�wH��+%W��P=��J�)FCWo{����q�Dm���]q7�������;
�K$��?߲ZӁ��)���/|��UnCf���E�o�S5@ԯ����yoǓN����Ù��U`��d�:5�?Z�R��e��j�ɎQ��û��~V��N)W�t���%4X2�2Q��æ/��N����F!z`H�7[h�m2��uQ��{q�c��w�;_�`:��"^�,G������Y�x��@m� �Y#��ZLII@�w�������:P�*��������T|C�9��7�+�Hf�&�zٳ�[Y*���wB5��>��<��Ot��}#���7�7r�O��[�L�ȶ
E�As~h�dT*G^���%�B�R�޼;�z�_o��r*�,�����	dMr,|qF�?�|��X�f~�7��L^re�<%\m��p��1ٚڢ�9��Z�t�Ќg�8�4����\�7�t"�h�}DL�:�_��.:c�Iɖ���.��:X�O
�̊98_��|3��1@7������N}yEj��?�#��sR %n���[0 �%"C4��Ѐ�m;��m W')�ɝj��~�i$��F"%k�Mὀ��М}��������p�ظw����G��<
��o�P�;�[(�i���Z�u�w l�>?�p}�ɛ�$OŔ��|ޱ�7)�2��~e)Q�3��HL
�x/*�fۣ�\H#ս�@TT�����j޲�S|�GPc<�� ��?`F������#��Ǻ`@�߫�܎���!)�v%r�5Q�o~4�yr	<��5��/�Ĭ���<��&/^7g�}	;��u����{_#���y,S
��S#��~Y�p�(�C0�yD�%�d�_�T�^��"��a��0�X	s��i�W�`��(��|=r�G�+m>���K��7���������׺��U�g�$�\=�j�%/�U[<��<O��P��B��NӴ<<�A�����U�L�.|��@���i�EH�ߣ*6��w�m+ow��Uw���l���>l�����Rc��C�Hge]Np���S)2#��SX;��ylz�_iq�>�01S-�H S�is�L?��W����.���}���ܡ�X���r�E������mT�'$���t,�������b�cIr��R8��-rJ3��3�ؔ'UN&��10Q0c#�2ߜ5�RL��8X`$�\Q�u#��ѴK�b���t���P?���!�=�YT�   ���~͞1��T1]xj�7�.� �|��J,:q����H����(����c@�j�)a���a��3>��t�a4�q2�ѭ�Ul����^��]c�]�5i���yC�
�/D��N[�@Z�^���0��'dϞ ��/z�3w��P���
���o[IE�]D�>ޟ�k/C?hz���KL�s�2�npe��l�|';F��޿ܒ_Ǝ>��{iM
 3��J��K�k���㭓;����'��Ȫ�)D�N��M@�Cu(^3�
��6�����|��q���)�a���}\��Uz����y�����_�[��,���Og���C��I����xg/���V^f��Y��Sݧ�Cv��Xv$���ӝ�6syt,a�ɰiC��r��ި��t�:�6����L��rV���R���+�=\ 
 3�$lN��0��I�P6)6��	�6c��}��1p.�ؑR���=�_Y��2R[����A��� ��n��qF�����~Vb(*v~���~����N�=�H=�ғk�$ʳ �=y  I_��S�=4t�� �u4�S�a�����ƒ�Rޥ�:�5�څ���MeG`뇢;��X�����ۭ�����[�/E1-�j�d�C<<�+8p���� t��Bݜ��,pi����s���#B5��yH�j˘��UD^jIF#"���}����+�Q��`#ѭ!�ejՄ�"�l,�Ъw�=7j����J�����4��X5[]�i݊��H(®�On���(�EhQ�B����O�t����P�p)���+��_%������ީX#�xq�����)o��Ҥ���8����k<�����	 �79��z��r����mh�T�V��kF\�zWڗ�d�P��Q,���5H)f3���%����	����*��{f��K�/v�a5p�7s}c����`��|[��ʞ��٩\�㹐�����p�	o~�{�uc�#�H�}��5'^�����7��-I�����$%�~^hT[\�88!AMW�?a�m+@0o�sTY���}�2�緁0��o�vT��T���%�#�d��, ��֩��M;���=ʯ����>Q~�QREރM�Z<�y[@�8�o��k���(u�	���ȏk NˀbY�F�;Sѿ�p��$JI{�0U�l(����Dai(�Ie�c�ٔ�u�<�%�΂KL�������Q���*�W7@PO��=DqVEs��W��������ϣ�k^?ۚϯd�t���@�V�}!C���CƉ���tB��1O0�/�]}�cz�b����_5z�h�z���U:�8�j/�}'GU�_�����}�Wn���4Sa�&I��d\�U�E^d]mwh����p�S.� �ȑM����{�H8"(8�&_0�6 ������L���T��A�%��ÂQY�u~lV�xF�\����V��Np߯��u9h�N�Y��B��r�`
h�9�3�#{�J�شૻ�e׷��ԜP������
Y�����G�y l�z2��EPBOB,ā��#i⬌;z̝�=���J��TV�:E
�R'_����;Cs]�|ޞ�'�qup�0B�x��[`.]���+(�H+�=m��:�;��� ����<[~1�#X~����o�H���F]��?7(����|k2�����!��J���@ZzU۷������{���{FI}�����gb�Ҧԩ+�(�Aw�M��: �X;�0}��$ϛ%��g����'X�d�"ad�Tv^��u�h�XJ�L>_'+��ٔ��B���5�ܽ��IJ�q���6A�}!ϼ5s=��H���Y�crs2#!�=Q�є�� 8�N��(��)B^��0.��\ev�{|B�ߛ�/T`\Xo=pm�\Zb2��I�V��B� ��ShԠ���P������u�,�O�c!�lÙ�o�$�qx�K�� Q��B�к�ܭ��jm�A�Cl+����]h�_���X�lCѥ�VmK7[�n5��?�[L�r�w�6���:TK���e��X�GBg�-�m��Fٌ��*TSfX. bXJZ��gl&�I.�ԝ�Xus��8ů�����VΞ��7H�l�GwǑk������5.P�ǉb�����>�g9���}W�a����y����ފ�h(�F��<i��!��*G�������K�s��x!�H����}��	`U����|����_�h��#���.��A��iq�i�%B�XN�ܐ�d`qƇx��Y�l6��-���o�)��� 1��`�k��@_���"q��<�U��	��������G]�I�,2�����'C�b�ǵN]U��DK�j�(�+��Bs�@���t2�Vv���c�iny�eK�ĢT��ODu~}_��ξ�y̋m;�6������3����|��� Q�S겙�J�N��h�u������������ʥ�>���9U����gc�&逾��4�,���Ϯ	v�{�+ϧ{l`��bL��|��v��y�4P���0�G<���d�3(J�%�c
�Ӻ�Zi�Y	� ��N�Ѳ�?����}�)8
8p���%Qj���G�j�{7R�_�u
WuR� ���y�]>:V0�d	"���e~qt?:�ׄ���X[b���l�$_{8�f�?�I��̩j��j�H�q��N����/t2��~�W��ñ��B���`��>�>�����Lz�ڐ8��to��b�;%�� ZJa7�)t*��A�_up�;�ňFV
��
:~�@���U���5����@̾�+Ds��H.ǌw�ɫ.0�jm^���	jef��v
�\�:�A�@�K>4y��0_X*��:��~u2P��v�oc���4�$��τ��T�Y��aWJ�*�hnG��13��,5v�]�G�ï��&��X�舅��T,�����~�����mx0��]����w�#PKġ^�>k��р��Sq����!W����֜Ҫ׈���dB���Ĩ�r��l�iA�=���g8*���ҒQ�<�Gy��LpZAEOGk-Ha��c���R��r+�'�s-�tX�}�G�Igky=�rt�C���pٖ�ҙ�*�t�9�$/�1���/�e�v��1�"̛�?b�26�5�u��A̪Ms��u�8���������lkV��	큪}��u;g��d0�q�@�(T�J��!�	��8� B��˼*�7h#\Q�� A_-��7�:6Ť_i�*�h&��,�G}g@�]Ğ=Q�x���i3�� �`r��� xXTN�F�>� ��zN�*֦��8�t(-5���!=/ �͠��a5}9ӯ@��z�����0�-5#(�ť�yJ[����#9:�L /\��%ܙ�Fi�{u��/S����4��C)R�16	lk�3@����ž
6Eڸ�Rh �3�B�����
�ڦ�=��ab�<�j_3�	��FFQ8E�/v͇f�+hh�e�R�JK��A;��a�5�䈧}��3&t�R��js�)���	�V��A�+�r.3v9�c�#̎^�� ��|]��$���J/��������u+�(}G�j��)^\��k�aO�H�s�x�4ֶx�i�Ѧ��_�%��!".�0��P~��Js�y�>�6�G�� R���SH�}�N�2<����R��I��#ZЛhТ�-�2�x_EJB���}bl�$�#��|ݔ�A;/,�͂�U�#Y��89=�؅KxF�T��#==��f��A� ������p:�.�yW�0ן��v��������C� ���Q]�)?|�u'�j"�e=��p�W�y�;�3�AD�_�)隨=]5d�9�s!�۰�J�EL�k���|�>�¸t�����)��ԕ�8A��0y�z����|�?ק�A�5~��G��T�4>�ˊ�_�N�!��
{A,�q� ��L�tA�0��4P\ZLݨ��|��~�Z���A�ޢ�uº��:��W�C8E��
j�A�y��D�š1��=o&�i+��5�-A�����S����n,VKe�z�_v�*
8�b�˂�4fe���?_��wҚmԖ`^tg�):��"���ּ��8��1��Z@�c裰�3����cBC�j1ϯ��c83��m�q��ww8�ŀ�(W'�8�Z��Z2w$�@�g�7]I��=�¢z)���#��~gF�~��8�A ��4�+���� B�GV�ӿ}(��D��'e��P�໴'$x"��hbC���',�q8��Db�:C+���fl�z	9���3�X��Å�BQ��0�u������u2|��|��i}:W��2Q���x ����%���2W����>sM@C<d��Q�~����g%͇+�9i)B���Lo��W+��\��T.�Ű�KfX��xC"��>�RƖ����5�����eu=����{ZT.�C����j,?ӫ@��&��ޔ
��g�j�]�(�mb,��!f}���&�Ȃc�o�V�R�7�Q�e�j3U����8���)}w ���ů/��V����\G�����6�Uv��r��^KV)B2�
���:ܩ��'*�Ç@�y�;c��.P�m,Ni���<�l��7i��k�VI��<��O�)�}�F��5��+ح�gP�_W�>��d�O �w�$(�3 SKH�*dZ�N�CJ
6��~b8a��׍���ˈF�1�Uf�;MP�J���g�����������?��x
u�!{-��k���O{nU(ɳt~a����PnIy �����e_s��T�Q��o	׸;���c�DCeZkO� F�	�F��H �x�qq��ʯ�9}.n��n}1֪L{���l��m;�˿q �l+���3����u�G&4��c�*{��˘�7w
!��Q��X���ji���6<ϽoD߱-y��;� ﭰ�_l�gm�#�2L{��z{�A�mf�&�9��*,:_�Ë���@���c���`Ug�Yj��|kO��}���V��hదuqtaĒ�-�l�)³n� ���"ȏA��<��a�%��T�0q��O�}K)Mڮ/X+n�����.�P!��&Ys�	����6��o�2*v>&%c��X�v����ꔜe�vq��bOJ�fz�ܱe7�-��R/���Y�����1�<� iY�%�*7T�4�p|�v�(B��m��3nL��D�������?�����`@�� -BH���� ��=����V��y���	ϲ�Ro��_~B�+��s�����BW�SZRA�G[Ρ�j�,&��Q�����|�_Hݳ&Y&E�t�Om� �Rt�F��������ms��B�&��0ܗ/O��l��O�.ݶQ|S^��|�t�3��6$i�T%��|i�O�Hs��EJl��@C���A�1
��l��B�Vޱ�_8т�0����X/V��I?��׿e�O�&8�W��^Ǽ�s���D�XQN�j���r�G�I:�6Xx���j����N�ЯN}&,�(+t׃p�nP�vZ���
����K������z�OZ��U��ֆSdKCq� N�_�1��q��ߨ,n;s^�F4����hN�
F`���lVa�x-��e�)4���e#��W��޹	�Kڪ$�!5l�j�������������j86�����
����ٯ-����6��~3������6b�%W�����@���u��@�O�:���ΦK�R@k����)�3'R_՛#B'4]�S�0��éV��_����I�B��=�D	`�t��6�R�>p�U]ǫM�lZJW�fޑ��`�EZja��c���x��C*lBáX}�q�0�* M��}潬H�P{!�+��%��6jw�z��u��wx&z��E��;�HI9'�oU��� V$e���P]��`�T��0Ҡ��7I$�
��J�Ǜ�3�*���=�G$��ۿ��
��v����,C�&|����P��DzoF��Z��Th�/�^����� r�%�LƵ�K(���l�#	�P�����΢��j�U�~ג`���В]u� ��1t���Vt�aP�2z��|V�+"�8�����	\�,�{���P�����;�24����u]ꆯtR�g@oAQ������l�)��i�A���I����lXJ1���U_�3��v���~��$Z�뀡��84�5��Z�,+7n��l�	6���Mh��=˃[�u�\x����0�c۶r��))<`-35I�j��8  l��������؎����1ɷ����h��(s�n���~�l�Z���6��+gN��V5W�ML�fek�섅���։;��:�M=�G�N�t���j�c��-:lK�k�2�����Eھ�v_��m	��I�6�뽨�1O�����+9�^|%#�W[z�Z�� o�ߥ�	� �G�95�����{bz��N�X������ꭆ�^9�ʟ�4Ź`��d��9X{��P��o1� ?W�ªO�M�1S�8�ZY0�Y��U���OO��G��e����A����*-�+�]Vz�|��EīӁ����\�z�3-�՘P����H�n�����Z�\��}y[�a�څş��,<Egn�;B����i�6�b�u���� o�2�fE?�����Мw�zB�Q<������;����F�[PM�k�~�ƈ������xr��}�B��[�v�%�r�/�[ �U
��lȪ)��U�p��f"D��8����q���pk�57�Q���Q��o�:{RC8z�#�'F��c��
׎N�J�� Ȉ��J�f<J��f�S
�*��\�In�k�	l�3��/��Jj�,�a�B���a��W�����\�h�4�H��ˮ5^��n���c1��2�����{&h뱩��'�0R��o���^��ʴ)f���>�1HV�,��Nx��;د��˺�� �6��z��U����*;ac.�Zn���W*CT���i;���gm���"GwV��ղ��l�%�y"���α�=��-C�p��g ��|�۲���^�F���������m�~zJGq�:ϫ��e������z�;������[s�u)�d�rh�>�%7H(m�%=�`��{�}s��橱[������L��L��b~��Q5�{~���I�O@E�#{�F+C���v�W(��e���4�����s��ڋu�/�⋄3������]a�/��o����1a���^L����\;�y#� �I�>g}EwN������68�l�7떣2��`��3"��Խ=~C\�I�01"� �#���]!IU�[�K"�s�֠80��)Z
�lM��a\���W�m�0'��8e6t�ũl-�7��t��ٞ�p�t�e>��<A@mX�!>)GD������>�R����.�a� G%��g����`N۩����C.�]Xp�|v��e0#���͛;L"��|^J���	��.}b�F	�e�d7qa�5�+�2	�b�C��6���%۵���D;e���8T0 ��-����I��xHEG��}�TB�B1�~-�����jҽ��C@��� > �t��$���1K��6�4ݩ�ٞT�������y��pk���bX"3z3,>V_:�4W,J���T"N��0��0C��iG)v����w����4"��5�*o��[����X;�)@h����Ds�@BjXt�X��.�B�H1�]�J96��ݜ��ʙH�g�p	�FP)|
ˈ�t���R8
f�\6EA(�w� �P��@i��	$�V˂��6��p�!?{O�j[<� ��Κ�_�_���5���%�����S�����+�_�U�B8j
�żP⌱}|�>6w2�,�����,M�8	�)�&��s��zc�jq(�dn9���g�@�x�i_t�R  ��1��A�� s��PJ��¯�%ao�5�&�χ@����v�!l���sl�]I�7h����~T?�\l �Tr��u]F��"7���}5)��_��_l#��̺>KX�]�����n[�,:gN$��#�uv�gW{��=��~ܠ��o/��m��9������hJ��#u ���Cg�ъ��Xl��rU`�(͓�#�O�iC?'(x}&��)~�����|Jlm@�_>�O�t=C�
p��y����h[��1˟�ͤd
D�D��Y���\<D�бV���8�#h?����R�'o����h�� ��������
���,���q�ɂ��Ծ�jF���Z/��9
�i��H�[�1�@������x�����(j�{�H���׳�\�w;q��_��؋Rf�d�_���Q`t��F�/�o�%��Y�M��?�����e�G�}]���4eL�!��w������hݓ�Y}���91��f�jgϦh��P�HF�����hX
�.���.�q��	]�{�P�%r�N��\i"G��	�yBm�y{�Q�QD�e�mݛTS�s(�Ƿ�W\3и���Z�G��C9qQ���{o�u�bG]5���b�M%#gad\_5������-�����W����b�a�cdn��[cV��פ��Z�6���a�z9,b���Ӱ�21�S!l���=���B`>��p�����/H|Δ��&�J��6#HR����Z;jrJ��Zb"����X�z7o ��+i�#��Ps�O�1�KW���z��Ւ�]t�88�~
L�a`o͂�WCoEOG��J	s]
{L���U��]O��4��+ t#��='�[ǩ
xT�@� 9L� �'���}��QLb����(�]kr.%�k��B]r�-J񚷦���[*�c^^�fx|�H�a
��z����FE���uo���@�-�B���6��Y}��q�/r$�@Uсd��o����9OW��8��ۿ4��<��߱jY��}(Ƚ� �^��+��Z-�9�0���&�����iP�1���C��q ���쓇Ye�E��C%k~SY=c����tҏ؋�-Ҽ��(�?v�r�I�� x���Wx ]�ө�l�����TKL��-8�jTN��_Ud�v�E��1��<�E�л��#x�Dn��QV�t�:�Ȭ�2��-� ��XlD}��4�a@�⢼8ޓ�1���_Z{3�qR��]�SsQlȼvޟ��V/띀��Ώ�'�ae�2�� ��(4�J�� 廲ڰ/�z�<��g�z�bj{a�Hh�Fο�c�+g���bi��A��}����6�E^eO�eJ!�m�Y(u`3��H��o���!e�L�YoejW(�&�}Tw�M>��#b<�Ɛ>�Q˨	��4�أ��vQưI�o���`N���H��� �d�S�<�h�w�S3%�T�FK�	��.}de�6��S$;�@�P�(��g`o��"�<)��7������ڝ��e>�6�^T��)�.\?�+�^�
HΏ�ǌp�
ޒ�½�g��X���c�dF:��қ��|���޷��Q�N������!qo?�/UQ�,�$�{�L�\��t�PEy�h�<�*�[@��z����aZ��g�k�ô����@�#4n'�G�T�����W�n�ft����� �h��\p�DJ���dJ���QUl�[�I� ��?{�-[�!-ȹ�_��o����c;����~]{1�N��ꯎ��bqLY�(l��1Kӕ�����������{��se�p4Vw�W�v��ff	Y�a�.�`*=y��|�K��ˮ��ţd�.l_M�P��i^�CHWH
�9�\{�٭�Pj���1�>i��(���Ġe�q��H:�o9�'�C����F�Ĩ�0�Ñz�njlt�����G��c��.��2�h��
1�X���r �S�RD�ё��i��9��:�Hݽ����O���C�Izk���u_10"3���Ӹ*�'$l�\�mM$S�g�|g|�O&�������^Zv�W"�����Ʋ:�	K��g�9H�K���x�Nn����D�MTM�R�ԵW��ځ��=x/�N��!}�jw�F�Y�5���wjn��oa�K�.;������%�Va��l#����1���J�6�4�ŧn�
���F�6�qe�/�8p:��1�[I��X]>5�9̙�:o`�?�q���Y�N��5���n��;��%bl���.{��j����Cc	$&��/�m�9���iQ�0:�[<���d�'��nTws7��#��kx��c�}{Ԛ�T�#�H
>x�|�"���ᘡZS6�z(*gX�i����N����v|���g���n�
<�2��q����M;b������pt�(N-�	a�sP�~փ&A4�~�����EG <��Wn��I)�6�Ã��f�!�����%�������{�9[��{ `RDL�G"l#�c;Ⱥ�#��p�!�Ϣ��,��z�W��Q��[Ӂ)ܟ�&��V�^?=`� ��b�xq��X��D�3O��7]lY�3|޽����B�MQRs`��� ���hB�G=9�(p{M)!̻�/� �ؤ���r�>�ωМ�ks?~�1�^H�Zc���Cj�&w9aW�ʷ�Ep Ӭ�q_����XK`�s�� �;H��KX�Ps?�޿yR�p��okm	Ɂ5��M��{"���j�X
2\;�v����5�rt@�h�V`��,Z�	>��CjL �����~����z��x�q����`  �ޥ{��,�$9)�Q��ڰ1B(��ٴ��0%|Ɔ�m��c�6��� i���_TFxÙ����\�9¦�� ѣ80?{?F��D���m 7	���܍�.����N�=�P�1��j�_��݁�Q8`���"x>_NM��ʃ��&32L/O�(^���`��R{3MWV�s�:�y	'��ٱ�6N۫c��ԝL8V���++�3���N�����Y�+��/���*�n�CM�,����t�~���!��N?)>�WJ�?�sP�~�N�Z���_��r�A�|�+=L�U�Zz��[�)�����QNu���v��ߔ6���da
X� �$��TU�yq�����b���~�.�%�9�i��1�6>�#l�8�*"���8�j0 �=3�qWQ�d4���V�U����!�7�L�7,�
�P�@�i����"w0���/_�1Y�oP�.��|�28�Il�l{���SfVF�[���ҏXv�dW3ݙ|�@�`|��'�����o}~����=v�=�� ƒ���q400~�@��K�Je�����z�IH���e�ȸ�����w��V�xCJ	9=����^�����W�!n��Z�b��2�D�.f�M{�R}ٯN�pU��g~�t�R(��.
��#�>���`A�^�)���B��	����@�B�
465H�����i�$��a++�Cn���dx�lHu	0� �T�?2%|'Cb��̨�@)�
��"[�r ��H�Vtg���)�%��B��X�Ub�񠚧&�ˬ�r�<��L����S��:���?	�R�[��V���4,/I7��vs���������<ha]����C����/j����������>-o�A�<�\$0M��i4XsM$J.?���_9��mae���H4cO� �����)�^Q�J�I؉p|ߙ^��^�_��3�S�`3�d� � �"��z� E��=\�;�v����t��ܮ��\I�A��{�������35%-6��m��e(r9F+��>�`e��������r���S����rCj�Į��y\��4�P���^}ι%�5�h�)C_�v�H����I���˶��lԧ����O�eCe}�	>��DV��'y@k��д�q�?4�Vz�n���<*d��������U��Q�&�d�
�.n�ޝF��8*K�U=Y�z��%�� +L�i�P�W��=��]�� Iv�]�o��,ӛ>-�wAp!x���!� �� o�[)�wB��Q~�\��{o�uF��p"��F�D�c�_���S4���R/�_��7���c�:S����)i�`��0�[�9�nJU�0�����?����!�3M�:�яFS;ٰIq������|����A� 
e�k��kq=l,s'��)|�T̈́>MU����EZ�~�sW��a�J���	�yxY3�*ρ�y
`�"��h)�D����1��!-��k��F�T����,YeU��p����p��H�ټ���C�Ր;.�o:��/�|�m�q��sgWMXV3��q��7w�����P�6�/#� �o���/��v�/PY�\h��qf�V������Hl�Ll(4:�[��W.ޑ[2�{̤���;�|ߏ6���ɛ�C+�Ex
i���s�y��p�� �,��ֈ|~J
H:�E
y��_cK'��%���|%E��ya^��4����ت9�F}A��}X��@]�b�]�ε+�W��9��~ 3�a�)~-Ɛ��O��U���܊��xL$h'|z�^�6�nľ�ZY���<���?��:���^�ӱ���m�L��B'm��H_�� ��4l��pW��$����GqLᐄ� ���,@s�6���>p�uƚV=�?�?���![��+�b�����w�^1��~�¼H����	���FU��]�p��3�t�
�?*SU��I��;�(t�+���@IŊ��0����/�k57�ɵs�i��D5s�z�q$�S7_��jS�&�O�EC��Nt"��
w��3	�����5��O�l�4����0�[I���I����7���=��z��R���h��<`���64	P�.��l�Z�4=�_9��r%���@B���)�t�����P��9�����n�P �1 ���sǧV��S3;�p�ocY:��)�]����ֳ�6FbB�J-+�:OK���"y�?�x}�����O˼�}C�Ɏb�4%>츹Hs��x��>��ۡ�3`x�w��;�B	~�E)�Ä���éz<Lv׼��P�,���f�o�s���Š�:g���ɼ��F�� J�wF�� �z�z��S�SiQAQ@�{*�!(���H�Ŷ��ȝ�Xಾc{.��
�k����Ԏe�˧�@t��lԢY�V�މ,��z��#{���O4uR�zr�%���H��6�eْk�#J:6��`Z�o�s�FhE�܅���D>��i�W,~!F��0اp�d��T����KT$���XL��3�W��t�i2�vX�>�n��M�?T����<��d�z����SX��4hk�:�Bu�1��{ޏ_5��� �������� �Z�?�s�T~����4�g
�;���8��w�/	���[� �.�/I�V�+uf�T����3F!���2A�����k�L��i.�Z{�UIu]��T�+��Lb�[�*�e�1�����[��@��s0eTDD��`6��o�O�g64��N������y��z�sڎ��r��"��ڻ�P�X��_<��מ���7{x��!�p�ޕⴇN�d�.`I�6"8L����)��F��C}�WTA>S �Y~�$�D�{(�Na�ןϮMw;
~��c�4���k���I�H�ܔ)+��km%=�z薜C9������N�uN��"0N���$-'_S�`K�}��ؐ�e��}�0�ҭH���&�� &r�.�M���!G�#��A��i�&��6/��l1D�l���w��ݘ=�K6�j��Z�Y�dL�Ecw��tU�WV̺�E0x�l9��D����;*U�������_M�.�p�m�ӌ�q`��A�vot��!�^��Y-�{N~@Y6��/�hp��C�za��_�s����L9���,�m�Z�}����Rj��ADTgJ7;'K�q_��Sc�?�*�Ʌ�'諛�i�z`��@� �-�����j�g�\�'9*7�![�����@eHX�җ4׺v�y�R3��羚uķf�u m��4eV��j	�g�����7����Y�s�Z���F�������·�`�~N�PƋ\���/�����,ysi��705�X��I��{z��;��;S������-���%}e�)�:O�tC瘑wӻ����	�ur��< )+1�_ǫ&��_ׅA*����(���4�	��Z0"�f��#`OL�U��ҒI�'-*P�h����	��Jh���;��?�e��G�B?��!��G���L�D/ȕ1�S0%fv����,�O/�5i��n�Br������>�����I	���3j-2�U��n$�Tp���&@yP���d:7$YΏ���˗�ܖ[����H+r9�9Ⱦ�M��j�6�d�+�~�z޷U5�S��$��dE�;��xH�(_�T,����Ḝ#~�)�ӧ��66���\�t}���0Րť�iG_|���ι��}B-B��k"9g���S�s,+D>砻d�\����o��3q�:�Z5������6L�q�� ݧEv¨�α�cVʐ+�0��aup�A��$�}�#�e����]�*��T���'2�j&�=��w��V��X�=$S��/ע��D`|rߟ�Dօ��X�y�J��a��_���o ��ֶD��r.'"R0}#?y��Q�ɗ�*��ƴ���<��'�fqI3d��m1Ŋ����� �!t��V�԰�䙓]�ެu�bLq`��~>�F�,�Я=8�Ug�S�Ҹ;);����sޑ�K��/qE(_��������.��]?�8�E@�$9���n��i2+�E�{R��Ao��ћ���P�ؐ�Z��B��HtAE�ޠ;�-_�;G8	��i��<t�u��	A��s��#�?��5�I�o!V�=�[$��ǿ�	��vf'��O����/���@��Rv��/h�HKѼ�v����Q*�Hǥ��4�طxI7��}�߫[c���Ƙ�jc댎��������<�sz��E���]��f
~�6�4�ǁ�QAK"7��*�t�<UG2�����F��!>Kw�3COyE;�"b�rF�Z@���������k�2�p������2&�,� 6�ܛjv����.?Tx���
�	)��(�S��_`�t�O�
�^�U�//:9}N	�Sr�ȡ�>�ܘ�'������6y��u�%U�X��^�M'�H��(:�4�$<2�ޣ�r�/"]�e��S@�πЕB�҇ĵ�\�E�
(�Y�F��%=Ƙ�mT� Y��qV�d�VY~2cS|p!pFW�Ԋ�%�"}��g���{V8 �:k6ps`��1�-�Ғ�,�n�^=�����K���\κ��b9_=w$���{�^s�&k�� �4�E���h ����/�f}#�~��T����n�>H�n��m{r5쀯X�ޢ(`T*��
	�wf�N�X�}[�]��bO;�8���DT����������^��d���ۭ]�^ze\�����4ե�I�ʆ�p��Ug#�cA�&���W��_s�#U,-��@�Q���22_J��͋�{�2�{Mo\�zJyC����p_���\�܃9��n����7�U��z�'Ǭ�6��M���1cƂ:=����\��<y�����h0�ƿ�=��G7��z$��}�y��eQdz�C��2�<7�in
��
�1;��%��BvRb�e�JA��FH��+/|�1�rJ��Ύk�g���3Nی.�F�w���'q3�J�h>�4�2o�,�<�=�z��
p��պ������v�!�D�(4����-����[-mf�h~w��&AufT�v[H :v.U.be�֫m�[4�)�M�:�v��	)�������nOR�a�N���ҩ}p�;�����Wl��qӂ�jn�8~5C��G��C�V�r�i����"S��ȧ|��6��y�z���_mR��I�m��n��r��e��U�n��#��5��y�a��Ǯ<hὡ=͸�yc�46�G1m5U1�_M���vI ��t�?�l��jӀ�����W�i���Qz�E=�8�#��.yR��Ҋ9Ew����Qd�V�F�pCm��''dHrQ%Ө�z�m��!W���E-oB^J�ZO�F��"��[�	�7����\�jfߤ�UI�I����\����I}hx|��L;�Ӈ�oc8�1�^�{�BL����7���V�n�%� }M�i�5��� ���hp�M��bB���>J��e/��V���"��j�Z�b�p�66T��nY�G�#
�H�[����p>��0����MX��Q0n�xD"Ć��O�sM� ɹ丽%^��i!=Í�O'�??�����c�W���s�e-8���̮n���b�$g��#�`�%�R6��JC���'
ӴXJ�c��(<��b�t�BC�˷�_(��谿qʸ�f}�db ��1Q��Sc�B^Q2f�6N�$��v<��uo�(��;��yݜ!Cʫ&5���[BS@s�9,�. <n�?$4{qzۂ�S�`�'k+[3w`��NpI�Y��k�vF����m5��Ax���q0����0�h�sf��f<��[]喍�gYC;_QNL�O�;���q�]0Wr�ܢ�g�LC��9w[x��w�s)�:y��o�0{�uIa��1����b�&��������'�Dؚ��!���H#�O[�����v)wqߺRO
/��7�v%��|X��F&�t�����A���:Я;�p�Y?F�$:A�8���'yx�����4b�DAW��n�	�5`;��KW��>��r�a)��@�;SF�	���$-���)W�o�]&N!HI¶�@�)���8��݇��4� ��TR"ʦ4�]7��%�.&�.��k^�:'G&�ُM��<�@��F?��2�_� ��@?��e;�L��O'�c��4 �樥eW�&�Ò����QNH�?<�+F��0�����)ּN(mۀ�(' ��Գ�\&��^��6/.f`��o����u�)?ceӑ��¶�"�!�O6�������J�8��H�ߏ瘥�ɫ��v��Ɗ@f���<Þ��k�"�W[X�B��3��}����g�C��q���1��{�uBP�͗�b܈ڻ������@�(<�x��>$����`�I�>���px���k�x��@4ن�ȥ���%��P���U��\!ύ/�9\d�T��2dx�5�g��l����F8d�O�!��|ł�>,�0��גV�������C�4���:;[A�A,�@�\U��!��+��,.|��;F4$��jP��Y�|4r��-�EK����(g쑬	��ş�����S�^�o�����x��o��_KH�^*�J;a-5�Ӯh��5y�ډ�{�{�8"V�5�+"Ʋ��e�]�.fd��rr�mȬ�I2d�o��u|��׬�>��M3��f�^M��� j:�+DF�16�#�G(�uN�m	�j�'�B�LY1
A�D�lkd��.-�&F&��X?��䪻)� ���xo���D���~��oTOUT��`tж�m'�!�HVqP��slJzS
�p��8+�+`<��?��vz��B��C"�MǂJ0pkRO�����ɫOϣ��|������9*G�8��Y:�U��-����Ҳ�u��:�>�#�P䲴�˹r(�]��%�"z�˳v&d�ܸ�n��d(Gᡗm@���b&ƚX<����RW҃jYa�X�G�����L������
T������T�}�K��z�l:}��he�зpg}v5�i�(�ۤ�h����ⰱ�}����#G%��Dg�i��pjC?�D��W#kv�LxJ<��S�Q�������P��@߀�Гu����_C<�YУ�w�5Jk_�zj��> �a��>��#|-�S��RR�3<�di��*B�.�hCm��	i�`=i�9��{�R`	���_/���V��z[]Q�Va��q1u��o����,B��/��S�c�D�Q��������ԉu����t��S<�0AN�Tqݰ���-ƨ��lPW�#DF�7�1��k��}Em��*�E[Q�y�3ȗ�٨�����;�€�{��	��(v�����~z�^D�����Q:�,�� ���B��d9��4F����dt9@m.U\�Rͯ�@�ܼ�N�0ºb� �z�X]�i����������z�b �L�����:&��c���!7_���7����Bi�"�"\Q�y��F��^j'����?��v�=- 	����f�I��k���YYd�#�)��д=:��]�"V譔�ZEg�%����*>�Y1L�%���-��uS�.���W7��?�B�i�v��@k%��gqw�e�
�W�Ô½|��b��2A�:0�o�3��/���c��C����>f���H҇[(1����Q�����٦B�.W���0kb��0E���m�����C#��7����g�6Ö
����5�n��z�s�ӛ5�u�Er�[�4�g�:�S$�g�x��ٙ��	)�f�����V4JAA*��m<��������h��mt2niH���U���yd`<�r�۾64FC(_j��鍏�ǰ�Jk-¬JW�L����0��+�9K4z1��>�P=�V�%�rh�:q�}{^l�Kp�+TOUjZ�nM��,�n��������wK�8��8��|5��t�N�@�]�q�cw���$]RO���8G;@�V��I�Y��oD��#��U$DS�GW�+�l9�.���o��pf ƿ�B-��U�(l�C��]"z�3�Nm�륰�G�� �@P�ʫ��s	���ܸ���8���s2�PlWqF���D^���R'W����Pd��c�o1C�A������.��?r7�ep�G�:��W�,�TW��r�R>M�4��KF٫���ػ���7��v%q[^��D�^<��� ���r�K��{���ş�{�<ZE�glh@$��}D����c�+]��-V�.��B%	��c�R��-c�#�zT4Q�E���o�6�<�q~�Oi���D��B����C�E����io�/��a�J-��+ώl��LY�����
�2�Orp/[D~�������(��5*vO_�7�i� B����1V}���ާu��2�F���5���6xG���-H�A%,Z����$@�{p�#��P��/�D�-�,��e5���������ѯ3�k�=�3����ɼ���`�Uz�肺X�IL��t��r��gk��I0��/��=B��&AJ/�V�~z	��xx�E������݁j�����C_vK"��@��u�=�����;�T����xU����kq�W�'�Lo��P;�Ε���,��T����Fc? 4�	մ&`'�����v%il�)��"	�5�TL,�|*���`�OJ�,^o�0GَwC�̍-qqXzh5��~P:�4�a��pI& �$)|0�g��U�:�
�A�~�;i Z��3�D~�e���g���X,Ϳ
�X|_������}�y��c+�R!0�P`�4fA��L���"�Xk�|���ư�5t�|��t��D��>�{�t�8�@;c��a3P�<bfᎃ!�U..��s���ߪ�C�֢g�?�ę'�+<��K���=��uI�]?K]^�^�g8��Y$�#Az���syk��)�&*rà�Q�2���2�Yo�߳�p.��NnA��؃�T�>>��W�}������u����� �β#�j�����������ě����6TJ'�w֦�x`�<{�s%53�Vo���`�G�=�J�n�un�io}.s=n�H��L��r���fX���\��}��kVX�j�B?��C��OK�����MH��'�NV�"y=���	J��vy��%\��7]�r�2J_��$9or���~�ޯ�\@Z�,���faH_U�z����z�/���Gy��6^_�!��-.'��'ɒ��W?|��ZR��Wm�CޟH������X�Y�/V$��A=���Ti�~�n�500�'� �e�J �Vޝ+HJ�C��k��M�R�K@6`�=v�R_;�<��3�f`�l��֟<��6(_�6�����-���p@Q�=�hr�K��Z7F�[{�-�슣�����ž��[:a����yv������yƫ��-H���M��at�!y������3�Fx#̈8mi�^\��onDp�ż$Wi8��P�?)E�"9�����rmv+�<A�b�4�����x\V
��1��#��4PRG���,����1^��A�]�M��`Zeb���}��!g��in
{��@���%�NAzIi���a�j,
�D���(XXd�Θ��53��35�ݮ��ӆ!<�O��܎2�������bdu�)�PY�~����l!������S��^p�X�;��� ��� uvG�����Y�ǊWޥ�b�Z�֛멻���5��8i��$�[���g2`��B��4���o:�C7����I��p[�k�Ȥ�	LА7:U�iHF����Rg[NX�:����98��ϐ����G��:-X���0�����V��I5��$2�
N�.�n��kק�%_C֤��]�����/S��Tl�7�ų2��Y����\زx�{6�2&&���`��U��4΃u�Č#�x�v����2�B6��o9{]S;��!��m�<����I���d��"XCk!d��P}�}�����#�nZ-xء� �<�6-N{��6����9�\�+WY���K&�t�����\�ZE0)�ؔE��
q*L����O1�-��։�u����\��hp�Ӈ���
)��D+�|@N��G/^-����C���w�L�V�ύf�c:<��)K���)6s:�견.�o9eY��p��Z,��b�I8�=���,\��#5z.��X���=�`W���q�m�o�����w	9��[�ؚ��84���D3��P4��d��G�]3�&�ˡ#��ֹ��P�Na����ǔ
���}C��/�'��-�(����bb:)����JНn��mw	s����/Zws�τq�N����ܙ�Ǟ�,�Ba(>|]�f����2��=� س���'Md܌��+!�$KԜ�=�y�%:Tk�m�G�_k��0{��́���ؒ�Z����RM�����X�~�������-�y[�y���ߐV�_�:�� ɭ�I�M��pA����.�A���>�����f�2g�ٷՠ\����{3c<�����f�$���Xx��� �~��$-^׏�'�h]�E�}����ǰ��>H<���EPĹB���2GW-�D�����u�k3�OI�}�L�o���ȑI
f���<Q#g�=>kXE�$.<TB6�K!��v	���`Cx�X�ոƟ�r�rf��U����N�q�����B�����d���<�cQѯ��Zi�~�NN��ɢ�
��&gfl;|c'�W����E���
�~�(���g��\GC2��;������A��f#E�~��<�R㨬��HNj��M�5�twGC�����֩�ay}7�i��s���[�ۘ�[�V`4�.'n>�|���F�=�oU�\�7�����N�槟���L��iwJ�~+�����U�Ppf�4����
���u�Kpm}OV�i��`�h���������U��l+$A����*a��#�]�^~�������Q�Ѧu��ϻ���W&����c��{9� �:/W��U�������_Դ���L�vQM)�%���A,c����i�>�����C�b!,:�NflJ�m#mub���o'�P�Ɋ���Yopg��]�ɌH��/	����Q}�� Kjf��*[��ȼ��p�D�7���W1��2X,��ȰK�{.�G�;��w~rW~6�ɭ�J�?�����������W�VpW�]�b���˞?�k�0������F
�z��xq���/;�Y�h�vl��1��5�c���eJ�R�6L?{�\����ݠ"�/�b>�Ǥ$^����M8yy�op�:�g�X�I�u�ĳvU�s�������MxI��ؗ�y�e��߼�F��[Q;
ay���1B�:���v|􎀹�� e�jiTN;G4���3���H��T�_��q����"�gE�b�5����WZ�[i╇���P�y*�@;�d��k����2��'�E���٣Tk	8��T��-���[�MuY��� fR�W�?�"FD Up���C�Ϧ��4�א;j�Y_M�x|�]�1�[�O�c��KD�"`Q��@�R�����)�B�1�E)��2Y�$���u�����y
kN����%�Դ��s�p���_]e�a�� J�Us&0�Ք}����Dĕ�\ ��(%)q|��*[�Ū! l-R��K������� �:�;ڑ�-?���8��4K��Qƪ��h}�_�^�X�3@'X��}/i��Dv'�J�N�� �g~7���� (�!���%8��Ho�ؤ��X��fo�>��~�F"��Z�Q&����:Q�uׅ��F����;�s���No��4��y�Ga���a�<3t΁��wF�X�T��y�cA�����.�Ѿ��9)MkĒ/�j��=�O�!��6�����b�O.-Z�t,�%5�$��i�Pő�,��kxig�uä�6�Ѽ�/��]E�4E��;7h��z;�>xq�ŦL3�x�Z�4,tZ!p�LSs��]	��rA	����\��G������緻�*��^��{|��ƽ�.���W�� �߆ٚ�<�eJ&�l�-����V�t�0B�'���Q�b~I�ʾ��X:ݐ�f�w�}��8�=S$�^�;���E��e��A��b��Xv�D�&���S4���]��S��`F�3�'���5d(@V������+�7�"͊����ÆX�"�F�ݷh�c�[n&t��-��N�|�I�K�-�'a���=� Fy�u�P/��X�`A���g��	#i��]�������R]��?]�I��(7q��B�PO��¤�G����*i�Og�/?St���� #�,�GPUsQ�M'{jc:��I�k�AH���͜�P��<OsחF*R����*���g,��P��)�����/�ꌧܢM��Pֵ�������jȊ�k���ϗ ��upaFM"�T����	KJ�V@E�y�V-U�H��S��"�^��2�q��+��!a��y���$��u#h��5���&�e9aM[J�i'�R�	l��{���v���h�!��`��"O��*96����6����B �ӫ���� ��cV�S-��` �gŅӃ0J�W�'F�rJqȣ�]�l��^9P�c��=��y�s�m����mЇ׿N�9	x�5������i6��~@���MdѾp-3�o�u�2f2�f�h����|�>��t���T1|H\��MΡ��p�Q.T�x��#�7_�z������������5�դĶ��a�	\�~��0�f�����k�b�2�]�Ҧ�${]i{�%�F�l�Dc;���zd���G��7�������UqeC�@㵞��j w	f�����V0�$�E|�*��b�]xՂ��dM��T^��7����e�t�p�K�Y4��!�;y���^D��	G��t0r	�?g$������1Q��st��[2Ŀ!]�Pp]�>�S$r�u��J(���L��C���<�����Wp�b\��Ǡ����W��A��T=# r��c+�-�H6 �����[���;���'�'�=0z������n��5����F�׺����@j�ۜ{\`��_Ϭ��Ϣ�o�3�yJ�ֈ����ά��W�!��{�Q]�_	�����+�{�}�-�:1_��`��j�ʩK�x`�<Þ
��T�,M_�K�\����A��~����=��dƑY�0��H��ܿ�Vgl��R ��:!�u�ҵB×�2�׀����]<�l��9�\��z�	���\��%�<���2_`x�4<�
!��}���qJI�>|��tu�<��뒔�p@�$Y��|.P��a�ϗ��X�OS1/yɬ�N�˻a��(7�zkF2WشA S،N�	���.Ț�rzZo'�x�x,*��7*'ː/y�DB����
x�������+�����$�-JJ|}�&{d���a��+�s�w�k�1���9ޏ��`m��%C��1��3�DK�1n����-��C0�V}7�d��hGj���Sƫ��9O���� ��g�DV� E7^f�Ǟ�~$h�G�p�A�^�0����SP�%�X���ג�^��.������D��fr~޻ �FԦ2u��p��}BZ��)>�-�8#�^7��W���2����P�h��5���,��,���	�Z�rԅ���j�}�G}�6GD |��e���!������aEA=�����7�1�[�iB!�Z�+)h���6a��}�T�vΐE����:�'���v��1 ���V�K��>/��z�(���P6aV2�ړ��4\�K%B��%>{6�� Y��g�Y�`]���T��k��w%���MإZ�T���k(w�]�bx-:���dD q�O��1�8̓*���T�V�:7�N����Z-�g�����AI��xP�g�k)w�Md0�d<�-ER�م�'���]�̞q]�l�6�JWg6	��cj����!F,��yN,�1�~����qxV�%�]�	��E8@t�&R�L���u�.4)��!DW4zY�Qf�^�ɕ��
7�k���ٝM"[�=3��>Հ�n��{�^��<\M�D��HV3�t<D��2� \DPV�35��St
+b�T��w������kֵ"��֕�~���,������o�b�< � ���t��)��%� �cb� }z��hw�p�Ƌy�ؔ|/��B���#t�ui��^���@��sp"�����˹y�p���m�	9jVU,:}#������/�:��y@��w�Ь$a��K�z������ZqNU��x�ls����=������72֔�SIA�>��f$��F���x�R� S�V���}AF+c�)����%��O�2i<x�d�*�*Bt%�ˇ��-�}q���n�0�������Ň[6���%'_���R���J�BҊ ۸V����NH��|��*n�;��(��0;��xZ��	^kPd�+JS������s�N�U���8�Qj �Q!'I���\Ķ�hy%��	���ﻕ�q���M+��v��Œ��Т�1���ԕ#�h5���j(~d<X����q�%	]*gh��⪴3L�쐠�K��1Br���D�y�T7n7���$�I�F��"��Z;�Oٴ�{/���~�m��J���R�D3-~n��׽�0�c��1d,�$"P]�T	���j1w�5��@MĈ5�Y J����oM���䎆Nt@y+_��ğ{�(:.0��ӷ�;\k�����?7�Ѻ�^�Q�>����f	��j�jtO�r�ʲFo�䯆�����cn@F�a�a�.�����00� ����G�Z���dT� G����KNsTEK���\Z}�|]�g(RZ�I�,�u�s�u(��)uC{C4o�H9,h����H�Áf�F��a�ͨ���.�[͠AsTN5��yߛ��WI�u&�"�{D֊%Hl�~�Fi��7�l��k���g��(�Con�U�W!"�̭'��(ӚJ��������^a��CmAR͔}!������ώ�7-g����.����Ю�Mr�
������C��Vv[ɐ5d���"��od�k5�<Ρ���K�C�&A�x|c��b����Ц��[֥E���ڃ��<��Y�\U����h��p�����<w��S���u�b�y��z=�tndm�P�֯6_�Y?췔|Ou¾ju�����w�%�v`yRS�Ylm����ga������ ��o�w�`}sr��h�.p�P&�/��@�W��O���eqC�qi���Ë��"��'�(����cm���|�%���r6�*n7=�6�eX��w����^
�r�Ć½�#/{�fQ�(�Gp [0ϧ`�_K�k�LDy���R*6K�w֋41��h�����_������ԝ�ɩM-Ӷ�a��l!���rd�2�C��O|��k�~��v7�G���&qXҗv�)���}ƯTv��q��A��(n�V�h�h��v���������)U�D��hY�63��j�?�l�r�b�B����1�9!�o� ֕5ԁ���@5;fvk��Vo놖�y�n&d��=�l��,�֘�a�h �c:!��,ɼ.�6_C�YuC��C��ٰg���5�!"sA��Vj_k���W��Yo ����.D��xK�,�פJ<���Q-��P?q�'D��q����1�~��B�,��I_�l̗C���̍hq���D]/�a�0�i�����@���m-}w6��]�����w��vc��v)N:�oō2_Om���NTT@`�1EZ��rVc�I1u|r��/
��7iE����<Xx�	"�p��:0�&A�u-��j��4,!���fN�p���LZ@`�l�J}7���c�D��C��*�ڍa[9�e�Z��A����/���!���? YC����)O���aV��S9m'�$��Ga��j�q3�l�z64_skj����υm�U�T�0�3�`$����ef�V�9zk��8U'l/�<w/&Nl<�S�^�3(MR���%��*���%��C�j��CI�����>�D�5T�-
*l�_��p��-!\��pQͨuKNqd��	���~�:��GC�,NM�7�����9H� �خ8��RP�ګ�t2a������fg9y�1f���pM�D�� 鶥Z/k�����9��'�� /�c�$M��Z�?t�["2'����[׃�+��%J��^}/���~ԵTL`-RK܍[+,���Fsx����v��L�Y�41����?|�Bu��B\�d�w��[D q8�MAxw��ߖ�9���NEs��xG�?�-�~;���k�dx<!��w��lJ6�zi$���R��'s<�$��TM��^8-�'���R���Oz�����m�1q=��T	:Ğ���-�5b�k�m�@���0G��B���'յ6O�z-��T��Ֆ�oT�o�W���E���L��Em]�?�D����@e�XS��ח��Z�U�zUnB��}0�p��HY����� �PVA�Bۑ(1�L�NGq��G~~���2MϘ���󧤑*.��Z'"�W�&�F��J�Y�t�{����A1ǻD��C#G<�~4[Zv�˜���Z�t���_ N_��3B9 uh�b�Fq�����:E/*Rkj�Ü<0�ףMW*��K��Tm�:�Մ���$f%7�g�-�M�jB琐{���eK~�PQX���V�V���'�̒�b�P#���G�E��\I��9��HfU�d��
B׾"�u�8��G���	M���g�L^%��2(�t����(��)����Z�]خ�C�7	 �!��Nd��tK�u}*�!�jF���j�
�	��=�q��rn1��`B��������$:��`����"��m�\=p��4�+������aӳ�s8eˆ��H�d��2��m1N�o��*Y�JF�ڎ*́j�{e���U���)4��D�F��3v�U�R�����bFX�H����~�)Y�� ���=yY�������Lڢ��Tf�"��G�,��cb�,t��k��;�����ŝy�ƥi���fު��*fg�z�9��@úZM����	n�ĵ3��z���86��b�^���:oX�n�� N��>�V+M�ѳ_��2�7��q��
B����(��u�؉W<������FR�-af猝�h�_���M�Wv�(NT�\�*��I³���"g�]�D]m����U6�	����E�x�'9V�EV�#�&itM�qh_��֓��	
�^��Lpw[�2��8i�e���N�<��`���I �si�$��YEO�"��3,��_"`�L�Ĳ+GA�E�Vt���{#Y֦P��#`��%mA׌�i���ǫ��#K�Wc���I��Ƙ�r{��2��j���X��zNU<]?F.� ��p�0Q*����=��`�*��h�m�y�J�I=���|Mo�k�Gd<���c;V�&g�č�.�lDU��PQY2aQE��x��3?Xo�?B��~?!/
����UJo�̃�;�J�'�i��(RLP��.��h���J}F��឵�b����
/Ě��١ץQ��*�y��`�)_�X'��?d[6��c11�������Q7��b�� �V�?����ȟ}���	y�@����A�H�I(/ �� �.iʥtw`�0���Flz8����k��>-�[ك�$8�^��Xw�o�I><��/�טzM=T�0�_Δ���?Uy1�",�?wm�t(L��;�B���9X�g�k��M�I��Ox3C�٢�GBg�nH��xO�;P�-�0���-�`詅}�`*�Ȁ�{�%��KtEz��_��>�� �j+s�QpX��3�{��MF��?ae���0�R��Gr��~	Z�r���fcmb"K>v��{�Y)��[ŗ�p�
.K�]E
�*y*"˷��Nȫ�,C��:���<F��:�}�}�e��^���]��=Ƨ��K�_�m�9�_��Zmrv�2���hyp�#���]��ͧ�ҧc͠5�X`��9�����2�f�xjXN\se��D�6ÿ�}�[��-����ͧ�a�$b�#�a������ mj��⮿�{�(5^VeD�C~�����49�\���]\�s$�a���Q+���^R����w�pv��N_�+�(��y������X)2M�0�ϗ ��[!+S���:�S�G��$�U�)���e�=����cM����`n�}�qdG'K�����#��8.y����yTY;�j�S��\�W$j��Is�8����������0������*��5�0�/�"��B����ҥ3�P�Ö�'>���+�1�`��a5��&��P��.���5 ��|�v7o+���Y�i� ;�p�>iR�n4�¶�ґ0�;BI��y��=�1DD��;�L��WY���C�)(���|��nc�<����c
�L�}���eh:��Y����;[�T@�*l�=/�)	���Q�!U\B%g�Qc���B�#�s�l�ܣ���Y|)ץ1RI{�Mܛ��O��@ n-��C	[@d�{#in0Az	q�3��������FU��W��J����mg��_fp��D�a?�EZU�F]�'X�E,����o�_��P$�w����D+��-��3���F���`�SU2�zj�k�ָK�d,5%��[R/o��ᘇ��]H�A�����c��W�u�"��Ŗ@dM��JJ8��ޫ��5���F��Z�(�K����C�O�y]���A�.IɺkL��{��JAR5����� Ueo$���|@(h�� �,쁒I8��2����R�U��_l�f>�T�;�+���Wg*���^�� ��8�H��6����JV���ݢkc�"YNƐV�3�W���ٱ�5���F.}���,����6�\�\�	)1+�-��&��(h��d���B3�����p�D��M�N�V���Α��Y+HDs���Y1V�ND��ڹ�,�U[��}d�dBM��0���mV�u��i�5-�-�3�d_d�,�.�?���0Z�h�c&�X�ʕ������0�		��"��8H4^֛���)�ke/ıx̑;��*��\�'�X���Ț�Z��+IX�q�߂!s���@t)�G^�.q�{�U��"�ʏ�t%�Ùm�Vh�o1����]`��6����S��~�[s���q�q�n�C����2�#$�U���2Q�l5msy�n�t ��=]=F�����)~��QN6>`6�F!�r�?H�P S���sV`�L��� w�U�(����qo!�`X��.7�8/�9`�-�\��8���/��,���aA׏#�f�G�hzHq�P�}��X�̑�Z��+��<���B!)�u���5��)�z�b���@�s����LJ�Om�S8�������ر]�Q�l�F�-R�a�[�����\�����sb�k �n��5������8�����DN���Y1���	N�T�+b�HB����rn�'D%� ����;�|�57�l��Z�����Q�]ܾ��	^du�8�*%:��9��<�fR?��X�V��}�~f�0��b�B��
p�R���)y5	�IX�q��u�Y3���k���9�!������9ԄH�r0σ�	�S�p�y���?�a|k��yK���]�`?����so�pp4td*| ��G(㾥u��!ǫWp@���{�T^��8�v�':V����/w�W�����,�z{��~��0
�a��5��D<VLeԨf-U����c�%0+0w(��ƴ�
| W(s�p�Z=�ޙ��/t$�آ����!|��Ag�Ѩ���}Q-�����E5oK+�������v`	�[w���]��L��@�K��:���l��yp�kD����}�;H�@7���e�{z�ܖ�"-v��֘��o�<`biR9H��\�?�)@�(6�= �m��c�c�C� <��4�5����fi���]^�=X|�P���v�F��j�Nb�'�1�H$YV��%���y�Ig��������7�g�}S�>�<��h9��K�0�p�����y<v����wH�J��Hhw��aa%������w�Q���o� �.�T�q]C[����!Dȉ�r��ae����hQ�u]��
d�~��},6ț�{prҖ2�;G���z/dM]Q8����)�D�c��6�l�׿MXƒ�Vxc��GU}X��DbW!��|6Z7|��IvЂ��I�8�_Wm�����u��N�>,;�.������ռBJ̪K�H�GA[G定�~��;#�
�Մ���$G+�Gt�M�;�y�������zq�2!��_����(�H36�ũ�Ȅ�UUS?�U�d �_�����s3�G�rE�D9=�j�)���fN��O� .��&�s�׵s������?�_OR��ԔgK�ퟯ��rZ�?�q�M��xZa"E�ȧx^0�@BV�ڹa7fY�xd��RL��u�{ٟ��u�J
 ��s�pKN�T��VT����p^��[��<��B$ID��ڕR�!��� �I�Í"���`]�b�	��'�����+DK@zZ�e;L$R��x�k�$��`��%x�DT����.+4�Cc��ի�T��]���>|�(�S5}w��^�ad���X�8�q�(�Ts�_�m.��%V�H��Y1,7�G0Fv_�۬�|=#xܔ��;h�0����1gX�=j"�*n�¢=�����G���|$<�tZ�n�T�y0oQ��a�.�/�4����"�!E�^ط��d�ŎC�V��Y��B�_�n$�Y��R";w��}�Z�I�}�sE(��?[W��=��ݜ+�/������X�^^_� �iV����5K���|u���/:]P#7�.u�,U�WnP��������D��E1A�i��*��AL��~6Y�R�9
��P�+�r4���~�J��%]G�� a_�B�-4L��(�`h������m�t�7i�d5�,��R��tV����t2~v߲�ȖF��_A�}`p!��R�D��}���2����]N�$#�q$U�>g�7ʰ�Ğ?�=���s��_?&�zn����x�	S�F=�7�;��*���Z,�چ��U��z��Y��6K!�x��<���T� ���j��h�9 Q*�R@��X���}V�*4c�����^��?�b �h��ۉ�,q%�i�B�o���Sr��=��*��:�aʪ�J����"z�;L��y ��:-_��5ݸ����w���ꘞI�(�P�O��7��)\J<Յ��?�+N�c�c��},���@k�^S]�c���P�����R����<n��>4�L0dmW�"z���?u����PfӨ�·�Ǩ�(�T�O������G�I������t�dF�)v
V�n���<�z� �6��D+�-'��6�%�
�����^�p�|>�wO�v�a���&�Q�@�(8H{�}'���FQ�.����,5 
�V���b�����;h�37���vs?�v���5�uLQ�)8"�^W30��{瞩�Ȝ�{�%��	�ώ6��w\���!�A���f��ˇk����SOf� ��B���x��ֶ�&��r�G�4
y�z�<�U(���9�
<��
$�D���_l�e�p�����Ց6���#@� �ӕ�]���}�(������4��+�Zo�b�4��n�6x�Z�u9���Bg�]�@��E������~Wj�ʸ�|��m8�!�~�C��j�7r<�󥓩s����x���g���Ǡ��xcM7����H�5ȁ���t�"j^��;��|������4����Cȸ��D��O�tA�(����0z���E�nDrP6������,�J��H�JFS������`�z{g%0�8�ؠ�}��ˬ�E/� M �^����j����ޑ
�_>(��cM|�r�j�c�LM�C��;j��s���3�r�RK���mv����{)Gg��z��v�Ա���lX.�˴׌�ӹ��)��R���M�`e���sM��k�q<�r��"X���B��������3�n�8����TN<P����Y��L�*׈ w��R�w�nu���՚©���������m�,��މ�z�#F'�r�̽��$	8�T�ȋC`i"���q���+L��O\�]K���9�5dzЎ�L�|r�������=ț�=�5�7�r���l�Q���ׯ�"[�;��%;;3Bl
�i�2R
GƫK9�d�f_h<�m�|7{1.Vu��Z����G^@���˓���f�1�p�<]'e��p������}G#9~9��p}�k�>�2uZ��jX�H��M�3�6G���Dͷ;�.��ыa���m�s��n�o�X�9h[�>	T�h�k�p�J$҇A����}K�����K�����8����lw��P�D��;c$z�Dή'v��if�O��I!SJ&�]�	�!yŷ::>
�!o�R=��Oߑ� &�����4��]{�i�|y�^a��.���d4�L�y K�j���&n�W�LEܯ)R�k��� �ߌ�E�d��x6ߤ-��W�T�ŻD�d5^֘Z�&��,��|����\�<Yݾj�#��ۀ��uH��lu�����Ğ��!,U�<���R��-k�G��B���)�5@sw��^��4��qJ`���1�",���.�,�g��?�ܾ D`��&ޒis��kHl ���<w/U%v�$U3}�P��9W7�̔�R��#>��	�äOrF�ko2���"�S���k����V�$0�^fz�m�@�ě��Z�.�63Ho�&z�f.Dcz���*�=�z��_�9�
۱�A
�U�AF��%�-;b�>��3֓[�S}�P_{E�Ld
���{�{�����P��J����A��<)�l������{������p��Nb$�?�|,��Ç�$�Nl>Ԝ��,�	�(��������>Ut��u��_��j�V-��������œ��E$sv)%�ZK�v��dצ��f���SPb�Z'˸���T(�O>���`���	�C�����!�l9�wv(�uL��c���mwuAz����Y��wZQ�oi~�M�}�k���@�Ua�0�/\s}���f���7�f{�2�4�z�;|0�C�A���'4Q����\����ݯW8�OC�����]&e	y]S�#o��#sv��u: ����u���U����Ee�,�k�[<�0T��Ʀ�;�3v+q��K�����An�i?��A�h�I�[]�^�4j��-�r�����$D���K#Ħ�0�N����UFh��kl��B�Չ��U�>�vV�V���-U{��n�b�w�N��a�Ⱥ��~��d�I�	H�q��c��W�:l�+}N���`��c=s�?��� M3�I��:�S�M��$(ax4)t���iYRB�����`�4dK����ᅉ��h��|���ۅ�Tj��_%��F�Pjﰊ0�
�d6�(2�ǱYr�r�I�����[�a8�/:��sӤk���6g�GF\�l�� 7��Ө�~/�����
�T�ik=R���e �/�kķad��x�ّؖI!Aƾ��_?R��@�(o����!�|e�S|����+��q��x�It0�����|e2��C4�gi��on.s�D�%��]�δ���w��4*\u�<��p�D�^�z|�P5>l���Mӡ����o3hʏ�0�B'Dnyj�c��^�V�c�0�/��#:�p����
��	��Z��.b��l��Ӵ��˯�����
�&�L�U��1���l(�[Ϲ!�	7��0&^6qiU�/�ɭN����A|2�@��9 ��\˔).=N�t�)�g)�}�R������f��i���6{�)F���	�q�\�6��.�4��&�P��Xh^�~>J�����u���7�}���>	 �z���8�Q�Ո<��f���[�^�j�)�1z������vZ
䱜�d�oD����;�ܔ۸~�K���PP<
Ծ�$��\$�^H�^#8Zm��H��/~�n�+������ೌ_s��Y���v��ʮL�j7f��V�Fi#*]kB��2��@�5�(�1%�gY�@�����0;͓�ג��v�ayC���60���˜!� ��Κ��S2ʅ�PKf�Z�ö��4B6M�����i�<K0��L౥��w����UNR<�K5��.����Nc&oV��r�Xk5u`����k�&r"��bq�-��1fT5vũ�pS��O��6&�~:�k��o7h]���[s&���n~���-�����_�}��u[��gIH��������u`���Ni'����1�h��z���p���a|��� ��P2&��Rb�SX�(�G.#��=�� �����|I_������,?P��2��S�C�<G�E b�`'A����U�C>Ч��i+p{(��Rw+�ɽ+~��R��o���W���M�T��6^��]AÚ~������8���um���)ƀ�v5���LC���ׁm5�����|�l̕��g�{�ƈ��k�7�r�,�?�,$���F���܅��U�3ˠ�;%�B����o�i�{�M\�ja��h����]�գ���V��N<C�a��3��,��5hx��M���ca@	��NZ�7����!�\��ki�	Z;x
��v{�N�py*yf=PQ��ɉ`�uW��ڱq쪪^�I|�@��l"�W�4��l��7��[��_=��HQ�OToF��򫣋��o��Dߥ�6(��k2�>O������G��r԰�Y�JE��{S	��L��\bA��[ǘgMu<��`bJ<[�Y���u�7�֛�$ZE8���O7�ޡ�*x�^Ȕ����j�[��71�z�Z�Xy�jr y���w@4�-"��LV�9R����.K7��ز>�N诫��`~9�^��୍*1�=B�5u��Mʨ��@�؏i
�Aõ�$�F�\�q��L���o��OK�O,'�͔ϭ@�5�0N~�Ԁ���f8�L�9�Tz���0�]ը�k
�U"��;_*�6&r�bx,Ө�0q&`J���RK�8,f��;��=�}����_��Z|j�O�E՟sx�Z����1Qc��K"�I9���'���� �Tѡ���B-v��,��L�9��0D�K����G����:Q^ݏφ�s#��f|E��C��~1@L��&{̷�����O�Po/��9<�*վn�|�ԲJ�נ.��.�����q>�o��?j^��k��ᙴ�	�1��`5��J��l�Bg�R7)I
��t�C��Xs��ꞑO��K �jb�%�P�d�9s���l��8������-���?�Bi��:7������s�H�$Ybi��&�'j��n��Z�����h�A�n�Þ
0ҷ�ɶ6}�� SM��X�����Ĳ�^�,�)�D4�t(�w20����������C�q��R�$�Z�n.p??/i	��:B)�����2��`H�`�U�i������Vڼ��W0���|��g/���M�z�f ק����c��<_࿱@�C@��<Fi��,Ge��G�y����m��v,���XIy攬��؇9c�9� �]䰝�d�M]5h��8
���aW��@G���bV��n�����Z�"�(�!�	���o���%��辨�n�E�mL�9G��*��l�12~�ח��7�붓��:ِKB�?\�O�����4��BnS(\�LQ��K:1p*՞�u����{ӻ�A�̌�#�s���r�����{/�]��έF�:���d\(B]�eVlǓ����
��x<��<&�q݃�&e����X��<"�_��J���B��h������y Uz���qz+��o���lUr8)i�ڭ+�����xD�)ͮf{���9&P�� WjK���.�D9�Q��Z�����N-}�u�|m�Hh�<X�5]�(`���N�4����?��s{߇���� B�c�������g�z�� 
�!0���_r�/��&B-��D�?�i��s��5��fc��i������|גL,aJsR���j���_
�5R�b�oI�
m�Q��6�v�0� GY^Z�ƞ��;�1U����۩�p�(M8?;�\^9���/LT.6�y����~��$"+7�?�7�Wg� *%%f�����νF~��aɨ�&��m}]��hH3��]����y9x���6�kW�"z���A8&E{�|�"ZDo�|��q��Y�rH�bP�ox=�yJ�v�w�J�	�%�uB�\ψlΔ�ǆeV5�Q[cJՌ�����@0;�����xu��j����B����O���J�5�x�����u��G� ��0�R�;�'�������N�x���zh�ǎ�F��
o@��������z6�*��_/������}�9�'1*�7�?&�RV� ��a�zu��_��x}N��E��q�Z�4޼�ݐ����>��C��v�}x�A��WC!W�Q�/�1ʯ.Ꝏ��R��5�G�2�Y�`�n�k+q�i�;.���V�����B�i��!�UT���د���7��t$�����f�7×�b-�ND�+P|�8�k[���lds��E"1�iSB��>Z�@�S>J*/t'�Ҿ��]j�a��@�w*����V�h�6��	D���?�"�Rbk���z@̲��)1t�qww7��=�r6p\	�LWw��rd������0�m�A���E��{�2�kBK|ɷ��ٌ݅�b?^`j�Ht�g��i�q��v��T�ųc��� á'6~"�P/�͕�+	��`�S+��ر]vQa���kMp��������Å��v_�_�
q�=N�� ˳��R��^�ʌ�� *�k�sU�MZ��``��7V׆"D�`�N�_Ş�ML�t�RpN��8�k��U��P���ɓ4���%�H�>KC��Ncx�{"A�>����H̀�rd�r�B����1j,	�9�ڙ�eu�_k\�Т�D)툶u�?'�[P�-��@Ғ�5�hМ�,�����?�C��r2 5V<�T���ګ����0̊�h����^�VujM��w�^���mDu{x�-���>|�y�I4�|�����糾w���]�.>�T��i8��Lh;�;,�y��� �E��+�4u(���q��U�eB�O�Bf�(��w٨�$`�U�-h���ΰ����R�DD汫�a��;u�U#��g8R�$�k���*,ل��S�8	E������(��p~�q�x�B�P<
'�WC�����U��.,��5U����?;f�9��SO�0K����>���B�\�X�4����Gj��`���~�؅���b5#X������+���z	���Jm�Yl�絲�{և_T
]`[/]�V�k�`���ʹ���;��U��Y�=%�D�����X��n�3R�A�����=e�{�4��@rz�u�,Y�8�mXMy�(��Br�r����F������G܊�w"+��t�߫����AY��X�[����K���mb����Vr��£K�dKk9B>��~��o�h�x\��8��#(��� ���"-Q�c�90M������]��$���!�Qe&w`1y��x.����a_[^z�/Z��aJ<�wq��)�c��N+i�Aׂi�,���f���v�v''�%��}PNO<�:��+0w������Ƥ�S#��Ewg��em�܋�n��}\w��C%�W�ʀޅ� -V	�0�l�B>�>��$���$��'���Aj�i����5��ěʮ=E��]��e���Jbv}�G"��Q���p��:�2���>�5���&�2֌��k���_Wn���!��PV�������ᄵ=mZ�|5%��n#k�(�A�h-TV{�C��Ih��ڝk�~LR���/�ʪ�e{ԃ�� �C�D8��%���?��S��y�fa:HM��?D+1��^5�!t��݃��&/�ˀ�����	Zq/�j�a��>|vp���� �J?w��;�T��,xh��Zd��ɰ ����EF���B�=�e3��X�>��H�'f�`Xg��&:@^����ԅ�0PJhbQ(䚶�9t�ko��'�r�Gn^� (R��B�sӸ��5�+�.�`C���}���Z� �����X���\a W��G�awiy�k��z�x�n<�q���0�T~��h�d��a_]�tBӸv��Y�"���zp^w�⯡��*>�l�up��M(��"]�T&�>a�p�/��nK]-�b>b�x�÷.��($�9�}�~:��|�zUW�a���kE!׀	Y7�wYc���gJ��[$^S.����<�7>�Og�M���2�e��f[�?C��=��Z��(q�j���0Ơ|�AN?c@��z�W��$���#����]y��YH�j%B���s;MaP�.������=d� �"|ِ)�S�z��(�1)���B�B.E2)7�%��g�ā��[�ӥ�4�l`��K�:q�mHb�j�X��x�<~^MK����#�&C�H�R��e(�dŅ @�A������!��S�LC7��r8�6� o��h0�&��� ��V#:K<��%	��0�r��A�ڹ��֣k�:fϦ�}X-�^�Ӆ?�dcC��]�)�����ρ7������;3>�ģǧ�]�w�F��T�S����c�˴��s��P֦�\�ݧ�o�H�L�rq�w�_U�$Z��bS{6��GO��&J6��양aݹ�FU���������`��Ws��+]W`}_���=﹑��EOLb[�F�ey��A��ɺ�L��5y2�	�F#�
XJ��G?n%Of�EE�C�,�va�n���U����?�p#�?��4��0ܣ<z��O\o+($˿��G�yi�S��폽r�[x��-Z㷀A���+A�N@��w�{����p��g��[vNh@�_�
pZ��y(�vW? _���}d���������k�<@6�_�5d�/eĸ�F���uW���g�ȃwF�����>0m�*1�@�lc���"�^]���Wx>�S1G��E�lK�P��4f: ��N�fqY 0���c$�vRB�S���Fэ����_"��
�YvyP��T�=��+�=|a���yk��<li� ��+h�( �JJ��<�1�P`���M_`x4;�j⇖��?_҂g���x1WAz�ޣ	fnx�8�(���̊z�H��C�@��9���jWE^���I� E#��T�e�Ti���|�NS#�vT�Ew��;�Uh�I�>IYAm.�'�[�cY�v�iEnFF�+V	;	��R���m��,�����_	%ȹB�a��T�U�u�Ds�υ�Ww���C��N�X� 	Y���g�O%ā�����ܐ�CCĻ/���.�K@��n�C��7�o=b�5QןM-�cȕL`*k Pyj�q�R4m7wK����^`�jk����C��m���q1�}k�L����A<^@�����P@Ԙ�"���\�c�j���X����a��rM���4�8�3���(S�������퀯iR�R��b��{UW�J�љJG�_[��gų��@\�K��Zb��"��VO��T�<�b��K�^�'/����@�&�+\��]"��F{����,�[��W"�5#b6(�}�T؀��[$(��'�;��A���3�:�m`V�A�kz\��@�����Q�|�$Y֙��88d赡z?����+�T�o��;��9�3���h�a�Wj Miv��6����iq���|7���[������↛w��I	�i����y3&o���e�!^���k�}�l~hT[	�BesS����w ��Ӧ�pN/�l����i��6a��m���5��֑�0�ۊ"Ď�F�	h��$�s��Ò��=v�Q�	�@w3�W�4���Q�ğ�L�6�ZAh�(�x%��U�t�ܕ����2c�i�����iL=g�NBn�8�}q�{��,#�<R�5�ٛ�Y]�kY�Y����;�����N�fT�D�w,�co���td0����u�P��P���7E׿x��εW���y�r� +������wMI�W��?	�v��}!O
<٫�S��'hlo�#6��e�k�m)o��#��}T�i'R�Y#G�t�߸(g(M-8�Q{(�|�PD���K3}�Y�Q�����]����N<��)f
����Yw��ݥLM]�~�� �&�*�	�VO��V�C�+.KyߍĉLi�5�ıp>���:p�²��8���O�,��Kg�'c�SrŲW�0t�n5*�]z�;}Avn�.������c���M:TRo("a�7/!|������&��@�����~F��[�u�4_o�_j��Ȃ�G~��
.�dIp�+�̢�{�9�t�2,����Ͳ#ڛ"��^��&M�z�^ P�UIF�a.��4o� kѽ��kzN�5tF�c�#Y.��~��ݚ]�WUo
L�
�!$���B��F�"!=Co��@6W���VVүJ},ץ��^u��?5B!�lƗîfp�:O�]&�����žB��=�����O��&z��_���2�j�u�X-�b�F��(�[��eS�uAJ��?�)�A��c&�Z�Z}��fQƵ �F��������z!q5©~@��P_�����^�\突�I�g��h��P=�w�M���ɢ��ȭtI:��c��NZ䭛���f0��~�_�����)&U�kPjJ��_;��R������D����x�d�]�f��gѬpKTsv��H�[L;4�J��T!�&I	�Rl~M�a�D�^�eX�3����#�,/��Rm��a���Z����سD��H6
�4���bX����jSy�չ=������s�@P�i�L��g־�.T�+��uōtu=S�!w�EڕMǘ����v\&q�;�Uc3�����y��A��ݲW��������݅B!�-/��ҋ�<ѭ��e��~d���%cb�D�����[M(�Wf�#쬧�p��0��NpjR&�����!�!�ۯsa���zM�W����vٴ��U�LF��	CsPo\�}�n
�Ih�x_�V���bD-Yr��~���σp�'��Y+&��Mװ��7р��� ��?aHJ�
�#�p���
�j�gR�pk��Eک�'uCE�_��.d̪�zN�JՈ��F��L1��p[F'd�v�n��o)KV{�1�G8�ϓ��p_Ժ��Bh�00%�UW!@�"��/�T����'�c�5g��u��0�.������n��@�JQ~�?�����3�Aޖ���S_i*���qj�b�۔a��ofwn�'�v�1�a1r��R��&���	���221w7n�S[�� O@eT,*����C�9&�Z/����� ӔW��<E�/D����e�*i���-B�73G%74o��uS�|�G:Qe%��%f�6QK��Қ�����@�PW1q���-��ro�|i�(�S�[y�W�\�%~�>�#�5]"�Pi����e?�� �_���2��戴62�K�����7��Ա��I7n����d�y���Ht�m-u�0r>E{��Z�.���������0=ٍ�����/~E){����GW���yϵ�9�K?�O�Ʃ��5!�
��E��yiI�u'��O_�B�Quu��}���WD�����4�Fߋ�W<�L$}��D߄�}�ǸC���>n#����E����N��/K"q)�&��v���z	�V��M#+�24����u�{m��?=eN��M�{c)��G�2��-"�����Q�9��o�z�k2{�G����E$���u"���J><aP� �n%ʶ�t�ɘ�˥��j媑UP�A�ݒ&2��U8q�g�YOXa�ι2�[���oĉ$*`���^�SAh��$4��#$�u6��(���R��I
���jŤ-�"h��5�.�g�aa0�9�^c�Xi�"�]��6W*@T�[(Z¢�ig�����u�a�`���X�v�^�����?�{�+�6��1�؎��ڽ��0�O�9�F�Σ��.�G�n⢮P�~�S���cy׬���#�⨢�ҧ;�K�P��f��r�,�Ԥ �ĤU�z�9���р����.�O�c?Y��h�#d"����:Yq��q�αQ*��i`�Cm��a��}))�BxFY��Y����('�6jO_�j�R-\�(�I���%ziN	�6��z�xH}�֓(y���pw�/��Z�ޟ��R�A��ѹy��_6��X^P���`�4��}���c��2�Q�[������F�R���B*b��D�}}��ə.���	��k�P�_�B�AD��(��6��Bs���C?L��*qP"I��ք��eT"��鶴֟�DI�����?T��a���8d�D:E^H���A��T�5�BB��@Y�8D�|[�F �*s�О�Nf�4i��%�= !gUt��^���L�r�v�/I�Ζ���6'�:�ٻ�����z�sLl�W�e�ws�]��t29�-�>����fk�x3�s��ͽKCkR-���H7C�b��e���S��c��� h�2�<����üQ��~�z�1�jV�KI�l!qrۨ��X��q�J����m���Z�aK���L��)e��ϛ6Wq�1kQ�}ucbob. ���Nv���%�J�>(8�壂:����^s�r���4���p��Ax08�(F���Ѹ������<����A1k�Kp�X����JLt��	��O�;���*>����þH��G�[ES��d ���)r&��Zi5#�j��o������R�b#I(�
��e@+�u�r�S�GƇ�������0����X+�K���Q"��K�[O�~��M&��[QZ������]-�e��5s%cMQ~,�hjA���%�=LW����D�7�C��J	��4��_͡�4BJ����/�0�J'ZFJj*qWF
���~E�W�6��!��yu�	�b�ۜ�Kܽ�Q7(9�+�x�mB�#�QpR(��@\`Ϫ��j�(�浠�
�2�D�}�R<�Ll��9[���9����^9�Y_\
�՘o8 ����V�7$1��p½X�F����z�\@���/��aC~iN!I�y�=���MGt�2��D�d��z�
Q��R���&�џ{Əq�R8+˙r�|�#q���o������Or0�� *h$q�8b�8�o���v+��?+̥m\��9�s�� ��C�9mڗr��XG�lD�\L�~� �?L���A�M4(78�ь;��)��\e�R�VW�\�k�W�wIDY���lgA%d�.�:�6+�g*�<�q�i Y~Z���?��Ӧg����F��u̓�!$C�ȯ�=���!���u���{�-�l,��C�(RE�.I��P|�i6������G�]�����iF>��z}��8Ӂ��u�O� ��0��	�V��nZ��F� �	�Yh� 1�`�"��bk��o������AJdLT�m;����h4կ��Hs#�b��pP�(_5.lxj�{S{�S�(�8o=ҟ׷h���Ē�����_zl.�?}o��ydƀ�
 �IK�~�cr_�v�H�\f"�����x��4~4-C��)f7!<�!���6i
�<�]9������~1ﰿ��6��&>�w�<Ol�I�b�{oe*���}o�� .������B���\wS���R�zQn���N;�6I�g�6�+�@j���5 b��>�?�\*:l&�C��+;C���s��d�0�4��9�
��>r��w�F�X:�xrwZ|�@�.��ne�-��:�;�zNl+46�,�bw(�����X)sǪZ��S�	_a�o��P;-������6qoU�t�DoD����b�_��[���-8����h���W��t�>0�t>B��*�d��^���1�D!��ͧ�J�I=)�W��֔pP`4���@z��g�i?Kयfi�ywL��t#��O�0�tX���£�3�':c�)!�Uԩ�$���{W�V��1��ed�Ծ'C�cN$��&PO���G;f�c#��b'Hc��%\�o�_C�4y�ևC����t/�ppDof�㧪z����0n+�R+R�L��1i3h
�;n'-��V���m�UU�bgGU� Oa����r �a�T�9� �U4����OjEޏ���߄or�a�m�U` �s8&�~���!ZAH��!B�:�n��ٴ(�o�3�}�����^��!eV�F�̡�2����K%�p�BR~(f�
)#��Nb�)(���0"[.
�Y6*^YM��5����@����q��E��q��{ǀ$F�����t2O�?��+�m�+��נJ[��qZ�c�!&�l�G����I��:��zf����/�DO�|�Fghp�H��2ښ���c,8��v�.N�dBOR�ir8��3!P��5\�ܐ�9���MHi|P	�Z����4r�����O3�p�s�9z�����%䏿B{��;H������A-^�D[˩�I��>,�r{���v�N?��+4��b�� ��s ��}��	�9vE�IQ�PBY� �[���r��0���qPh^�\���q|T`������B�
��,��`D
�zZ���83�̥�{]��}� �	~R/L���~V�Ƭ?�j��g�>Ϟ[=��%��*��]'1���^A�g���	d��@	a��<zI��!��~���o(d�C���m�[c�:�$�9>d����_��!��~1��/����Qo�F@�\�Oh�700ټ-Ce�*�k��Baސ����ʞ�A�q�n o��{�]lZ�����
F���k�J�'XC�PR.�:S2I&�[�⶧y^��KP� �*���J�ӥ8`����:%�lʠɻ��.8�F^��6�1�_����XS������H���'�{]���(
�|,f���:� R(���rEMh�4�H2�^���d��կ�%%"}�& �����|�v���{�]g���ȳx&���jxh5�C���E�ߝ�+�0�li����wQ9�E�B���`��N����[�N��)5ʍ�=���s�x��>�p�zc���]�����/��j��_�ݮ6����S(��O"aد22ص�B�aVqo�@ ���q�h���c%Y�\����%�Ɓ�}��%��+u/ k�f��J$h��ۄ�)5���jjIg�O�A�pٹ��L&:�R�e�]	���9t�k��e�N����+v'Е�$��jz����y`r�Ky�?�Wi���lEk�N����Z���ޢ/�NH��>�ղ�j���K�H,�Q C��`�[1E���(�#-V�z�x��9Hx��&�;�goy��:���퀮��bC	�|rF=Џ	O�}�X1��G�w4`M3XQՃ�^>����PKޮKU^I��������Z-[w�s"��/<�Y ���}�]ī�7��Sn������υ��	�4�CXI*�X��F7��"�qJX�2'�	lB�(?&A��p��"n�������9^8߻Y3P���fr�n��°�b�J��z��(7���]P�C�P�ٖ��P�k�+��e2�5ֱ��i1GJM��$ ?��]��.�|ڛÀ�����$K�������Fs�,Ӝ�2�n�������5�s��R��eD����}�}S��1O��"���=>Z�+���/KU�R)�y�����X>D�0�<����*������oevb��7!�&'���5����E���6q�*H���s_L���� 0	���@���s^|lY�!�����oS��5�W��Qj�g�_�*/��1�9�� 	�U��B�����n�t�U���ljaZ39bb������<�vx\�V�R����ϭ���G6�o��0畘������Mj�B��B���S��m(D�U\�89�L�������Ed�����<�A�F*�)��=ji���n~g��YN���$���'<&���|��D)8�b�&��\��+���7-��8K:�㠽�b�,4�(�Y�l�S��2FM�n��߸8$��2u�O�ϟ4��䦑�SsKrR~��3����&��=���13�:U���9��.2��2_����C�X����<l��9a��垝�g-��VO��N�}Ӝ�p��c1ފqk��9��SC5ʝ'o�	>웷\h`1d]�R�Ɠ<����]"(�u�^O�!P����e�Ӣv��R�-�yA��~��hqF�5ۃk���ſ6PN �az�����o�{zm!�
.���:a�&�%�g����L�1��ĈQ�n�Gu�������iQN�k������Tr���ˤ��3Q�#��	&��j�$r�β;��)���#��.�����[����L��� ��
.l�m�L{	/�Z3-GՃ���J�P������#��[�Ӭ\��������<�.����Xo���0�}\�
�x�~9�	��#��V�p�Кq=o�F�B.�ƶ��q��n��`o~SJ,z�P:b�j��7I���dl�Wv�PG��n���J�V\){����ۀ����c��8��� >^d��yvG\��F�����6��� �u�=o�/ �]r��G�P?2��e�;Z~���}�/������ �k�F��^]~ޣ��Ww����-�	�D�p�?�l�sE����~��V!�?�t,w�z-�_Z��՚2��B�}X!u� E�pe������d��G�u�����09�>L@#��A�[C�_Z�}F>�-�v>*��{�g���R��Z�o9���	J�=Q2^֛��tI����?T7�WaS���E>�C.�Q%��-35��iê�g4��3���8�gtsV����Ruu���K���f&�:fF!��t�L]v�B��2��38�������ӽ��`z��W��|�#���>���MJ�`��ވ�P�l*�����>C5Y�3v����G"3.
�k��2��Jl��ud�0��Y1Sϗd����O�%�Y�?A^DX]X5�gNI	m�Em�����0=�G�3YX�=�U$�ј!�7�;��"BYO>�l�C��b�I�Y�����/[�[Ծ/�j��=ҥ2�C��S�v��C��^ܓ�V	؈dه�����! =B�C��b�$�nI��r�>��>gU��p�#�LͦT��)�tB�A����cD?��:Z̠�RՋV�5��p��G.=�:�4 ���O$�� >����3R�t	��Si��2vx��ĩNl�T}�QM�=�`z>	��tơ"�ݑf��(�-yME�VH�F��:�K��B�)?����;"�q�!��2.���E�T�4 �_�#�K+D�}�5ܡX5
`9:M��������s��������??�/�s#��PDR��H<���t�:�����E兎M�"ѮMZv����%�&|U�\�W�%Gw;
uI0Y��`o#���6�Q�^�6Ԡ�-6�e�4�U	X�+`�P<=R4b�����S�`ڨ��<��˚B�r�D��������7;�w�Vt�vV���K ��,p$k;��2�(����4P%R��e�X���{:�t[�F��Wɐv�6K���� �
����G�ȦsqM�:䋋V��m q��y�����m�I8�O.�<u�XJ q�@����u[N�7�m�{lA QT;�*o|�^��i;ۏO�%ŗ�ҍ�;*�̊�,�,�&�eR���)?T�p��>q�J�'OU�'�b�s>Uz����-�Ɏ`=V&tLÒ�1��Ak�hB8�s¸(W����%Q����"�a��:��0|��_��B�B�Q4���CG�� #3h�G���rr�J1Ex���p��¡�]#2�wY�zD���|��0��^y`��]6l���jc���]�2CIL�H��/���Y"��v�hu�?�h��o�{ �t_���
K(���=��z�6t���'����Z��wm�*����m%9�{�����b/y�+�}Qq��]�}L��3���T����[#^�	U	�e��yN��Y�Y.m�?m��$[��;7�$��.rM�M���HB�,-��&#~J�!�`���S���wJUZ�5���UpZ��8�:-B�^"�=mw����:���W=_��^�
uZ��
Ǣ-�e��d��v4�|�4���+���ӜVgmYW,�b��z�(-��<�Ν��Ul��%68�Q�|{�u����O�N_��\�ʭ�Ȣ�D�0�}���p9܂A�:Ň�+�q`�0bP�)��e���������'0�����=�p�s��T;�"]��V�*���re�_��i
��ȿ���iă�:C�;��Qת.�}�j��aY��H�-&d��ܭ������8!�k�"�G=�nlx_GE^$�z�/��E�=5ə0@L5
r�w�Pv/�����Q�E���t��qfܑ�O����D��<���Wg��D�{����H>?��U��EHA��&d�	��]���Y@�r��T'������[���A����H�Q�zeEw��c5Hʹ3��.�98��{�R#��@��7�5��}����©�W�줼��	D�p���8<��ofR�G5/Re�d���]z`%�S�E	���j+�������O�00����8�
soQ� �<��{���u���� �o��ܕ-ʭ�-��{��F���q�:+9���E~S(~J��`���;#�3su��pF��o��iCݍ��6��uib���C���B:���W���J/	����25b����^1�`���5�,�'N��64N�#óN��;���Ah���zC=��:�+��"n❁���i�ͼ��������(�6��3�lD�fk�`;��Z��߫�q�tgD
��TN8�цt�x��%���P [7M�߲؄��&��s�/�*���,�g����W�h�O�xaf%ـ��e��>,h�$F����	���$e:ەm�O�K��R�����Md�n+1��%E����&$Q_�z΍ޙ��]��΢��Q�;�C�f~&;I,���@�Kf������E����e����:+�9��n�Lj��`H�vl�H��T#q�j��YL���t��nB�:�=T������b���bȜ��z&hp�����A���}?(�cP��1�7��C�������ɴ9�@�Q��f�j���z��EVӏ���oU�g�A_b�U�WC���>'63~)��Ym
��L��"J��E߂j6��{��뎠��K�[gfc�b��i���yĄ�Ĩ�T[Sl��<:0�l��v��&�X	=bc�ᒢ�5��Q�Vx1�dU�����Js�oE9(@�dj���1Lj��*�@}�xaeI�6��C@״*��A��5.�RS���~~tZ@����M����bzbO3Eb�&��1 _B���GEAO<���&JԴ�r7���6�U��n�t��Sh�X:鈈��fg��(�F��&�g�'	�p�/<����C����D��������n�eo��-5.$S�Q�n��M������y<~����Z4���L�m��,�es���S�+a�]�<��J��Q�'��r�O��ꅒʇ�N���a�mY�mBL��u �ʹp��ISueb�_�����1ϻ�J��%�X�
MҘ�n@����dݯٖu�S(u�+�dAr�쪿�!̪��W{������*�����ė#����we�Q=}B�6Rc��\,�@� -5�k��@�nkA�2G3|S%Og�8��e�eʛ��qgQ��e�N�'���^O�S�kੌ\��	a#�m3�	��SS�d�C%�mRo9����bo��,H��Ufi�j�$l!�u�Z�C6x8�=6ゎ\�f��^X ,�T���SEΫ,M�l���G�1��P�(�G_����A!����J�I���ͮR=6�2��;���H�w-��o��_��&ӧ%�9N�X�6C�O�<o��,�E�;�/g2����?���uzb��:�ȈP\�+4���\�1D�.����_k����"v�u`�L .����lVB9-؉!XEC*s�];e��y&A�o��vPhV$p!U�p޸�t� ���lǢ�%/����dm�죪{������WS���J�u��#���M�L#Dj(r2_h��<�N�MˏH�h��>�I=\�c�Pe��E�X���n�2ؕ��T�<��2�W����L��U�/b�PKYX{H����b�Z|?O|Ia�m{�M �S5������+*���� N�aP�A�;�5IJZt��D��eM_��+�ڃ�@�v&[�k2gۢ�'��G__4���Y|�����OX[R~��	��$r����%�j���@�+�L���Pgd0M3�=x��
G솰��H�8̏l�?�M�?���z��,��t�� z�E�0SM	2o���^9��'�se�<A�-���d�7Y4��Ѹ���FGA��쓠�_�Y$@u���r����ܐWJ³e�isv��$
o4~'I(�Xm��?oA��{��U�w���T�"c�fQ�4i��2%�\t��z�N����F^w�V[N�$���QV��sܹ$��M��͟/}=:�h�uYW����RC�*��^דR��|4�D2|��¤��Q��9>"��-���[�����J�'sN���5�5�� su����YL�a�W���� 3G�_X�&��c�,�ނ������|ԶM���������{��t76�����#�L�>톩C����E1m�y�Na0�xMn����m���:�%�C���mC$����I�u/�\T��ۚ�'(?������In���4Zk��5�u9�3-)��/{����dP�8�����ͼ��Y׉(��=B�Sf������6���=��Q��2Pi)�2����Sm4�rD�/d��r�/������t��ܠ�/�1�91��9N���f�ot%���ñ�/0aCӐ�!��k2y.YZ��He���W�^��(�q���W��x�R')�3(��%�h��u�	�ɧ�F��L]
�{���&4�$+�[A%>����D?����zަ�
�~^�����q�X
=M��G�7|�P���!n��c�t�"CԞ��Ҭ?��C����H�Y�Y�4	���(��>W0 �=8�M�4�iy���S. +�UR�g@�(���'�6�\�ωoS(��X�D�NHf�>+t$���0p��[V?z�v�3����J�=҃,������Q����*�͚Y�[�����H�8n'�熾B��!P̆ܼ��{��?Sb�j�r��5Z�_�mT~��?]|J�X�|Ӄ_�*�5���(�!�*]wP�Ua�P^i-�Y:�����=����`���!����Btx �r)0.��������*�{�cS�P�5m]�I�O:�%��)�H�}E�SW[����'{Tv��&~�Y���3;g�|���ZF�E����U��\�0,C�N�7Dq%eE�aƪe��ud��^V
):��嬜��&��d�-�4|���|����=R}�	�G~#��׽!��4��>�X�fSu������r�s�?�Rp�����ߤjv	�WFz#�*�����-���،���ߥ�c��	����8��iJ�]327T��Y�M���T\�e�偗1����MУ��yⱅ,�	�� �n�Q�F)G�1�<�p�5M��ߢ�E������=���A�V��q��i6�-�I)z���ƨ!�Q�YM�~.J�O��|�Ņ }�C�?�+ٿ�l�L%>'b�,ӽ�L1��h�l�W��U�� J����AZQ��Μet|sb�š2��c�w��q<�=s��wdc颲8�q�Y��YG��=ɍ8,Gl@pl�L��y�!�p�
N�]��q��l*��c[���>�2��p1i�3z�����r����&����NJٴ4D�&�L���˒Rͮ�\&f����V�����[Zs� �C��G�G�����$�W���)!-�eD���)�&�P�_J�e�����E�=Z�?���G<y�eUP��WzM�4DXW�뺻�V9�h3�iߧ�D��l~TWo>{�P�@��Sm6F�ʗ ��ig`o�� W�>f��]9R��$�IA�~6�O,��V}��7Kf߷FuU�PE~ح�K�%^��D�+
!��ɀ1��H��0��<D.�2���0k ;0���?���g7�(�k,����LG����~�Rа�{_���D�GT������n���Y@�4�e/�e�P�AD��<��\�٩��Nݖ�g��iV�w<T�?�U@?�ml��g��i�LtIkoLr*/�Z O;Cd�Lf� 1ܴc���	da�;�S��#rڄ����u�<��πx�3cN���ݷ�A��m8l���Y�t ��}�ϠE
I�F��J-ࠌA��M�� ����3�KxeO]����t�d�r�U��Z<WڥǞk����ݴOĨc �JRS�J��i��I?Of� �A�^����e�Q��ἢ�u��{�v���ۤ���P�GO�uqi��b3cp�����N�F&����X��OM˅��t�,'5M�ץ�4L�Rt�7�3k����(	�g2�.�¼KXɚ��gE��v��~�y�!���6��/�@��2T��ee�+�G\�]ᵑK[����}����(`M�8�(Ԕ�.�#�8 >���oǮ�*��,|�g���]�lyr��_�]4|�Ҳ���^CgK	�\;P\*w2-^T>O紉��kj1H�&�O�32��|��x����<�G�ů�/�3uO.�r^,x�>���p��|Y~��brR�9uV��[�D9i��12�
��(�s��m_NX�Iؠ�tm$�DT�+�0Z7�ߦB�1��y>�ʾ������"Jz�*����[A���f?��+�g�c]?la@UX�Z�K�r`�������L����D"&Y!�hV�=�%2S�DiYL,�C\e|��n�-{<�L�E�'����J!�Kz�V��*�����K;�WLd:���1�5�-0W�Б���r�4O؀m�D1���vTp���O���⚱��/�L��kq̋��cq��7���k�r��ӱ�U䩩x�����*���v�����u�H��-��-nV��X��=�>��;���]���{!2��ő.+I��S!��#h��V&[�N��X��ܚ��,��S]qԻ�Kpb���>I��ә��2

�3��/��]U�9ş9T�P���J-�юW5��Z�����)<��^�������$v�=U���TZ����[�*Q�Vv��E
-�?�K9՘�PN|�.���	f��-�ɤ;�������}z&����>�$�u��&���y��1�ǓM{Y߸��3��Wc擄T��6�7TS���Y~�IBN� g��a;H˪=������W��T�?'��Ǽ|ed|'�9-�y0/_F�7/ɞ�~��S�VK
�M{�������{���=v�j?#�+��%q�Y�P��>	>���F�(�8��"�g�P	Ŭa/B� �d����⛘�joٞ�Z<����#L(%9��m�}I�hg���[��.��@��`UZX��o`cl��h�e�k�V�ux6o��Īv.}*�v$ήܘ#�L�Uky���� �TO�}���hbk�U�c�{Q�Z
���}S�֊�i�p�_������T�Q�0H����O����I�}cٙ��f���1cI��,���Z�M���,�������FR�c�\		��d
O�������GY1���G�mk��-N�`�� =9W�ÕR�C���臖M���V���)�O�.$S/����8`�k=�����[Ox��_m�J��`N(f�ثzL���?�֮�a"��U/֎3�o�)cT9䫉U��o��	tK�'c2�i������)�==Z�F��|C��B���O�m�j��{2�5Vc���紭X$��s��#ߙ>��ƾ��w�б��Ɯ.��0h)�1�5��������
t��t�j]�Za�r#�VU���Ot;��pa������ً�բ��s�A}�S�,x�vI�<���[����c<y$��*a ��2yf��Y�"6Y.V��Ķ�r���T��!n^<!9�e*�gW�����ȶw1��͸5����.��i��_�� �f(�yY�[B�j0;d?��|Kf���S`�9 *(Q,C��=�bhF�B����^�܄#˗p��y�X�v��b����]�T�H�䴾��HX�KU-�.�����i�KB�~��rq�r��G�Y*�uf�A:ج�:�J���O��QK �< GI��.�T*.��C$D��u[z�
ŵ�K��v�U����>/�t��R�*u�B4zBR�M����~�����m�	�ǿ��dc�=��WgF��oȚ�NЩh�{��������Q�d�=s8���tX�;�>�.�u�M��:JH���
~o�d6���U��
B��u��M��N��o�c)9ϵ�Ug+���O�*�ġ��V��AbZr��u�djk<u:�d%~wq��#I�半t��C�6HBR�z�!�a�iN���_����B�t�a�jE4*���0��М%$�����3��b�<r��>�����I��M1�L0Z,�`+��&�����0|�I�EQ��j��eΕ��pJ��d�e�	h�y�����9瓰vH"��f�@�L�6���LB�$ +��8���c���wL�����O�'��
5~N/��0e۵Y��	�x~�Cy:v�������l[�~C�"�O�n��x-�|�t�GX��_"��_W��]���SH���(�ײZ���|����[�?�+��E]��ȕr(~A�X�Yx%|b���c&|��
�u�6�V�R�~?��LS���.uS7.Q������� �SZ�|�mKX<W$P\]�����h፮&O4t!�~����#P��� �2iGN�Ҕ5�����Y��t)�]�Mڰ�2��qӖ�KC0��Cj�p�|-�)�s�N�x�C�a�}�;��3
�,F����bV����,$�([�[���v��Q�Z��*>��)�v8�7T(1��n������A�x��#�S�I}%���Ӝ�[b�o�`%Ϊ�p}�1��r-�⏗F<&�L�~�	
�M<�e��ᄵ�X
\]!~r�,�4����"���-�p;��g�JԱ5��ۛn�Wj���Y�v��ߖ����
�hp.U6,�MA�Wv�Ҡˍ����)�4�fB"TWѧ��6���~��j��7.����/��ث.�t��	�H3�?�8�9P�St�z^D�z�F����'�v%~&ŉ�|v�	:m9���\$�z\��-�j.��%�	��%��{�p�Y���X��j�\�2�EZ�},�4-q
t�}�Q�'�us�u�a�����O�� �o(�~)/���}����%o�3�C��\��9о4eYC����! �b��f��9Tޠ`O��lL�G���'t�g�G�����m��5�L��V�"�p���/�����DI�u�e#XΜ~1��쿎xR�y�M�,��Iʺ}̓u��l��{�{��)2��7��T��H_0�C��P�����/�ߍ�Fr(���'ZSU4�$�u g_S����C㼾��@�H?g�m�z�$`����,�()��{�L���8�,��D�tz�W���`H�X�;(�5�饟6�HLJ]DmI
b�Y:Y����T1iE?vY6Ӵ ��N9�=��8	QU�������+٬E�zY%���k,����bO�2M"Ѧ@}��J%"��� �[A|༗ �%�N��`��d����~ȩ�ߥd����{i-i�c�i�d��~��t�溭{�R��gL��/:���h��$�$�d�)�S�LW����l�A�xB�C�.M8�"��ܐ���F�9�&����}�����B���tS\ڹ�V ���6����E�
&o*���r�1�ު+ޟLg!�rp�|���߫^��;�J9Gn>�61�	I�,=Q{���M�b�I�>&n��[�ہ9��:yƏ�V2k�@d#,�[f����q�x���C	S��f���*5z֜ 6��٥�c��c�aW����0�[7��hz�P�o$8��l��4h�g~�]&3��=�`��3�_wR\3�N��mƛ35�V����8	Z�P|#���%A�f�������Ajm�@�[��
ڲ�5fA�VR:�	� ��@��g| ����q��J�{�`�yg�}j��cf��Ч%����j�h��zeI/F9��a4<��2��?�3�O]5�bg0����v�q�{V�~�~��� )�(�Uȳ�;�2�ѧUW�a�8���]v��a/lƁMT�z&��	�S��+�5�J6�[�$�~�z6�)>�jԱ�i����'J�tc�8��cI�%A�|KID�(+���z^����w��'�`v�W�b؉y�2/b�p1�7]� �9�0�6��U9d�/�P���,I-͗-D8�x�8��S���X:��JHf�urr��&¹��g���E�\N%���e���L��)�����T��Y��Yք�Ocoim�ki [i�cm�K-בkx�ᰟ"����˒��%C����ԁ���X�\3�b�.�}�3����s������>j����Ȃ��;?C��@��q5�IϨIG�]�#�k�gd� ���_���c�1�/�痧�1��be���s���~�y�m|�>�}TT� P�f�f���ˌ#ϩ}�@�Yl���X+	us��7��q��Bq�k���Z?2�h,c�������{�kߧP�+i�<���5)�lɼ�:?du��F��͜׫V�Ef=�l^DřL�!��g=�V��#>�tV�*'���Ѡz�>PWK�S��٠U��>��`�p���>pW�݃Z������ L
�
<B�20h�����g��C�rn��3��6�.N5�T�Z�w�p���/Bv����%�w�v��׬D�^��0�X0�%P\
��>�p4�MDqj$,^dF�(����4#��q@U{P��5L���Y0��Շ��J,qMqeb��$��G����3��0�yԛa�M��b�ш&M�wh��.�h,�����_��j�:	0�<���+�����F�N'�a%4K�6�,�K�^���U�����Z���r^o��=Te��Yi挫��L� ������~�_�Nl��t�*���d}�1x��Քwj�N�G򮱃Hӵ�U w9T�@z���	��)$lݷ�c�|`�1�
��ٯ�����!�&8�,��qՍ�63����M����x����FE�r���UԊ�f[�5�"?I��tBO��g��f`��-y�XP�E)M�u�p�� [t���:�M���{ǜ��IP��r[Dy��`�Bo}��(���-a���-g-T�v_o=�9"��uVV�h�?ŗ�V)�� S�sb�Iu��VK��%��ZWQ��)�h��ޛg�F��n>�A��`�p�#o�~�?�l>��@!�&�`��J�����,ؙ��Ϛ����Y��HdF���]wT��p�)A՗�5y�Vh�f��[Qw�{�3�؃��(�{π��r��ٌ�$O/��Q����_���^<�d�Mh��΄�)q_����\�hH��^Y+mi8���&�4m'&N��D��<�h�t���b����R�ὄ\+u���G�|n���.lZ�Bc�5���n�?;���o|QC?�}w�	�Q W�њ8R7�cY��F��ňl��H �o�[�s���^�1a��glE�k�F�۶��"w6�G��Wz3�`s��E������$al�L��E���o�����Q2f^5�B�!�P���&�S��(И?MN?��
4��ّ�+$��-)ꖕ��)�!K
����`�R�)G���`�n: ���.�v��T}�J@��ɦ�1��hO�5��X� ����ث7?���x�O����B��+ o��	"��6J�C>)J&��:�T�C�OmK4��3o��^�7(�{ą�J\E�/򜺽��.��?�)���z��b(N 5ܱ&��|;<�����G��Df���Wy���m9��Ô>�7��&��ǥ�����ra'��0�]&[Q��I���S^J�6��Ԣ3l'��o��Y	`�����(r��}W1̛��3"�v��(������l"O(CR%��o�i�K
A�N�֔+��۫D���F�a���
���Ye��Q [�ae��4X$W`m��p��P�А.C�W���K��1ؾ�p+ȊF�X�f��N��ػ<ޑv��px)��[��L ���7�`�FG�ˆun�M�<��d���<�E�Eu����1���sO�=ZlT�A��FNPc�O��y��^ D������9���w�Z���(�B5�9;N~��>�ժ�2��������8�-@�:u���+��vj�4�c6��
��B�(����n��ݙͰS�1g~]��F<�������=�P������k|.�NE��>����މ��j�mV���I˪�,�7廅� <sP������)Fuj$�.�����A/�aW�C	T���o�Fct~K�>��-b��;��N�F2���F���5�/�]R�P�������"�b���>MX6D�+�f����'�r��'���}`�]��4�`���6`�@�I���'�'!��e���ռ�[���W|A��w�
U������s����9Q�Se�t�9��.U��8ۓ�f;I��c.<'^R����K)�)t�ܹ�ڕ':sT�`]�>�(����WP���}�n7����E ��bݷw�������z����[�{{]�fM�_����fO��Hm��;�j}������|���~�v������؈�UVq�n3���p�����̝A�+�6�
�*�.C���m�z��=i�{�毎��'/x��ΰU�[b�6	W��>eA1d�����$P:��wu��]YD�е/������*�Z�Nb��/�\����]�Ua[�ݖd��(�O���ܶ���P�5t�/�stN�Ԣ 9��a�R�1�-5���X��9m����=��m����T�:�^]����1�-U�\��R9b_����ư�6av��H(���~�[NA���`�m�+��OLU~��[Z�w��.��� �֋AOVre#C͢�{%0��p� _�q�PM�0ݪ�S�3��߆}�M�G#9�|�&�m��]�O��"��w3��o�6���s'o+�Am���8A�8OJTƫ�� �)��}\���ϖOl���e�����+�k3���L�,�m�r�	,U�{D}m*(�-O�vL��<��6B-!s��X�
kX�X�w`�!�$
��ܔXN��G�q�Њc�ڹ�u?�q��0@/<iD���{rUSPu�+z�u�V8_����f֦�
�R���4�J�\͕Ԕ@@�}��������t<�+��m��,~��N���t�}-�r3"eKf�.v��kFB���X��8���G�D�5t&�YU�x�F�)�G,]�Q:-��fOS/��]sz!z���jp �HA`�6#:����
��a�\ϐ���ɗ��%z �][BvB��%
��@df�Gt��؁ͫ)$�m7f��R:�Y�Rd���yp�O�q�&,��=��E���k!bQ`�,��θ�5&��X���Pyqp!V�9�m�$�D�/
��-��o�q�Q���G/J|�L�jf�a%�ҳ�M�LC�j!J>K�:F3�	�%��h��Y���~&�t�
V�Dv�X�A���(���8p����?a�ut��_���!�m王�-���89�����uy�m��z�N�I++o�1���3��]\U���IGV��(�!R�Aƅ
Z�AˣX''<�e
R�eԦ���RY�� ���4���r�`��W�/���G��8������c�4}֩:�NC����S�k���4��nj������פȆXZ<f��d�_M�L�`_+��I��.B1N���+3WB���{/�������y�  ����}Ƭ��#��Fz�����Ŧ���@�A������ �%㍗_n�z��Y����4T����ù��=�J�0 ��s1�G�>)��x*��;[�&����ۂ�MO���(`7�	���}�;(Ծ$c�J_m'�AL)��������*t݁�=i�Mͺ/�ᎽE'Ͷѐ]!�Pc�����65Lt���"�z��&�T��n+P@�[̗j�d��6
�n+ņ���$C��Ow)*��wG����#�����YS���T�D�l4��*A��K�BZI�GFM}�� �����Q�ӡq9�����w/���H���gD���c1�Fl��h�F��&~c3���:��P�z�M����R���l�(�Կ���<v�]T�Y3}1ʴ��iҝ����H��o�h�bi>˾��3BT�mF[�pP�4Z���g�.��6�"��Z���Py�����a�{����N��N_�}�a���M4��2��X�� ��i�M�
��@Pt�z�4�����:^m���G������Y5{,z���<yY�;�P�zO��i7�&k��(�QŤ2ŔoIX���z~�r,�V+մ��Gn,W��8��>�'#;u�b^��vE�����1�H��{Ԫ:�ћ��OI���B�h��Ҥ���*
$;�0_��g��+Qޤ+�"k���z.}9���\7��	;��%�v\d��|'uΥ�"�H�S�5=�{��>�o�1���@��}�O�"}o�~�YD�8�W�5K�6���;�a6"�g��K�b���6�?D|��¼���S*��YbttW��-v�:�N<A�|���J�1mlG0�Be�K	�&A��"L@��/����s)_����U
:yY��'�Kf`/_O�3�I�B�&����J}��U��wE-�W �����qpY_K��3�g�����B\d��s�lКS3�/�i��ab5"E?`%;wi�;!�*&�c9ިA�Z��PA�w^��1
Oi۠z�S;��xf%�r+[b7.�Ls_��'��f���a|�i�7�;dɶT��O��$+$�+�팺�����%A"�>xxLn��|��02 �TEs�>z"�Ӿd�զ���O_�85��0���y��Gw)�PC~?����c����d���ـ��p�/3�*MZ�:s�����z_	������Yb^�0��M���ό�r�e��|l��b�)�ғ�mY�wǓ�ei�i���zf`F	\y�, �دV�Jy�(�/�o,k��?�������G�� 1AQ���ҕ��X���>�_��t��-���Y����To��l�~���~��?��/�x�)�Y�[���!��BS��tmE^�q䜸�,^5�渉�1�WW�0���ddN1#��(��g*8L���٢�\	s~���9���Đ�=Uc�-6��[u����δ�C�ރo�>-q����!��^s̿�/1�����g�c���c�:�YFߍ��IX��#�r]�*X�8��n�$�_�2�m����,�Z��E_&��I�+u�2�0���	T��1��R����Y8�5�<���<Gy��K#7Й�o��k��х|ȸ�} T��q��@�]~iߖ��޸�к3�_�H�
|݋� u��fo�ؠ�W[ŭ�����J2��ߝ|�-)�A��t�j3�w�]���î�?��Kz��/�G4�*�D+�s�a]3_��yH�ܟn�����,㸠e �����]�R�fqb�PFY��r?����3�v�z�;�%r�O�:��nN����L�o%���U�����$ڌ�	���0.C6��+gi�R�JiE��{��y�1�J����Qrl����#��ƃ5߫Pz�҂O�L����g�xu������#����4VIU�MC �	�������r �RM�eN`�w�����\��b��×���l��*GF�"��7�#���7w<��{�b�J&
!*�K���c�6�=�\�P�UR�k�?���n�;���Jt��b��](M@�R)\j~3%�f����X�d�����G��|8��F+�����Gt3�v�Դ�~'�N��ǭ���<����Q#��>�@���s�S{����k�ހ��^�P̊5^��rX3.ѱ���N��qݩ����T8yv0-:Ub)��nD�j:��斢��5J�����#����.�m�0�:�ڭ�<�g`�T�I���KyZ��eٳ%FO�D��X>�WW�:$T�G��ܗ�����]K�`����Ù}ŋy4%��p�Y����|�����lÜO~�T-M:2�y��#�Q�tg��1��2.�MLc�8�|0�+i��f�r'&���P�7�~�U}ذ��1������'�a�uֵ�\��!Z@)�Z`��C�����:e��]��؞w�=e�������D�Z�d�y��}��E��rX�
���MI�4[�u�5�(��rR;�c��_t�zDX7؉V�<A�7���]��|�n��*<��q�1���]�8�(V6��0�.������Gq�?�$�PZ�O$����9���
�p9�
Qe(��z!�����q��#G ��M�� <\l(Z���eey�*T�Y��A��7�H!3���a�%X�H)vк��2�4����.J�����bh��xb�����,���r��[�[L���_�����ǳ�ښٵ�xng�;���� �%���9��	/��L�5�4P	��+�%e�w�RX��g�����>C�;(עÈ�}s�H̷:�{_W��w&���+�O��i���\T	*���V�v:�*^+Z4��VqL1ŻVzc�}�Y��>K��Ľ���X��z�5����*F�1b�\'2E�k��µt�3.�-�[�	��lKV�L6h�7}L��Y*mk �;��X��˵�B��8�����c'��*gI|��S����'����P	�гx*:�6�܆��~�nH��90����B}DwR��xq��8�������@�Q�j\�c��v���	{ܦ]ib��M[Qa����� >�����S���x�A����܃��5H����Y�£�R�?R`���N����>�
�
�t��@d�M��*&�S�����c���G����ɫv)��>l3Z�h�Q?C�h_��u�u��+$��[X�}�({o��2bw�z���e�z=�0K>i=�,΂dN�RЄ-a��/�a�]�ƬCZ��NWp)Aw�31B����>*+[R�z������fj���YC0<".�e�-��-C�̧�����u���3\k:�KM�=p��}���� \�<�����ZC���3�L;�}/��G�"��j��R���d���#�!��b[��c<~F���� q���T�\&I>�������
�^*+I�Q���S$��u#����gqL4v7��m� mf)��5��7*��=���s1xv_��*���k>鮤� [8v�s"n�#�d\ ��z���a->��/qu�	 �rVM�ަ/0#"��/���'����zȷH��I*���"M��3�����ٛ>�T�[�����@mo�S�7�ǕA��L�aR�����@80��y���@9Eҥ��s� �l+��#���{�2���'�h�1/�Ƈ��K����;���g�1��'(���$�l�4�x�qE8�D�~Â���y 9v�?R��gB8E�> #_�O�u�J]�h����ǆ�0��*俆�V���Kl?�%\_xY��/��r�f<�v�yVpR�V�0^��7/����@���S��2�����mr.x�Te��	��ب�ꃳ��%��&��yd^�,��Sohp����"r��a�HAK�_�n5�t�T��I�zNs	�U�����)����,��[�Wk��"0s�}�/��m�����e���9�MҼ��7�� ��Ƈ1rBEL�ԍdb�>��1|%G^M1��e�qb�H�B:ۤEN�,r�2���ꊆ�=�\ԗM�$�D4V-�)�|�8���i�v�Q�L_}������k��XX�KG�nY���.o�	]#)"�4"���P��G�:KD�c�|��1�U���=�9<�G��@C��-Y�pD�<Pĩ�xΓ{���{���`���R	�WCu߽?s�_lY����?�d�{�eۉ^��BxN��ՠ�]���@�hxx��G@�����1�q����.�O9՟
o�m󡭮�=�b�*.�h�J�]�ߍʥ_:xc���H�h�2�ә�i��dJ�ǝ��l�`pԄz�YݩN�<��p�YW�k�ƓvRu��U8 4+��#�������;�牀�S�s��c0�L��_A7���_00֌*��*pj}�ビ*�0�������^X���MSq���J�����8aR��$Ƅ)��]O�S�C�'$�=/�J�ͭ��3�����h�QKVHC�
A��^�3��t�B�N���8��A�^+��/۲x��O"N:�H�q�uH��Z~"���l�Go�CkIJ�r�MY����?�yVGm���n�EA�"����ܟl��t�Z�V<�F��@uk{*7w�XnhĐ�ux�^�	�t�S6{�d�<:�6������!s�1 >?��l�8���Y����͍m���)+l:Ϛ MĎ�UaNSq.�i�6QX	�#��N�EZ�����ҏ��q�V~�;k"��5�W�LK���)�`v)^$��^�Ƒ�í�+�	�A�g4e!��R��7#�+h,e��&�߿�插�1�/���`z:C5P��H��Wl���Pp'�;�Ȏ�ie�`�'5a�Z��M� N}��z���R�Z�9���tV��.j��n h]��̐	 ?��\��H�Q��}�m���=�ZZʙ�|�*I�TNl��Ζ�[�K�}�i�TՍ0�����w��w�S\K�)���Q�ٍ���]yJKB+��+��W҆y��׼#�B��ur��w�X��H��R��e|�C����v�5��
b��ބ�x������%��߯>���w�`Rn�-TE1@�T�F4P��&�#bzvݮ%M���S�G��TX�+�	�t�3�`4�&�(aE���k��!�E��q��*K</�u�J^����2BU
��p��T!�f��`]!m�g���|�X�t�����?�j�;Ϊ	���4�t����O&��fES��(�:$r�H�=���w7�Il�ڳ}�Jq���H��ʵ�]�s�$C�T*X�+�{�g����$��`3@� ������n�R��_�Z��|�fn�?�#,P��C��� �U&ffB���E#"� ˉ�\��A�=8Vm�}� a�G�f�}�������I{�e)��X%��K������ÎI�E�I��ލ���v�ө������-�{�D�͊A�p��i"h?�r���_=��9G��f�SG	͸�}���řn�a��g7҄���M����c)���e������U꤆ތ����7^��v�"0�:M�����bF5-��H~Kf\p�@�	Z���3V'@��3���<�᠐���]��d�$F�*uì�)�;��(�������9�C���#:d44[�/9��W�<<�Ɠy+Ց��ʏ1�]`=]T{gd�rD����2,�A�.ʺ�IQ-��5�?X?ۛf@�Aԫܴؘ�u�x�č&���Z����^������b��ʰ��9</t�9��l\�ژ��pK�����U��W�Y�ǳ�QǀÏ#��]]7C�&,�y*V��v��z�S��}!A�}�t���#Ddژ��4�-��9f���hI�-�?�J�k���y�-ui����6�\AY�X��i��
�Q0��
�!���8�T0��4Cf|):y�S�k�>	#�	��]�g�*�P�_�6�
Q��S�y��f��'������(*��_��L��9s�)���G�"^à�J5s��Ғ��{�O=AˎOa���Y��e��x��A� �#�Tּ�� �3��NJ�B�C󲚖�I�z���BW�T),v��:.�.5wX�*!�t�cZX�0,4�֠
�%۷#FS�xr��O���-�I�56
?i-~���\�ο�X�<�K��/�X�o�6�y���V9Eմ�>����>��NHut���3��r�X��G-�y"ąю����T3���}-÷ES����㤘�<q5E������������T�K����՝S�9�����nm���<���Y��F��[��S�	��ǹ@�N��5[\bd�cg��#����T�9����;��V����w�r�$k��x�����ą��ʱ��xL��%�f?� �@��9�1�K�V�Y����}�3`���H@ɺmW"��G����W]�@ӪwdE�"K�њ���K������'��y��9�Z�ӹ;�������
HR5�z0�Jf?j� ��\�e�R�����s��U�WQ3`���V�G�)����B-�/p�{�o<�M�-˩�I��1�~nL��H����ϽQJ�]Q�2_��w����퐿Ż7G�yi�=#/�����Ō�hL�2(��|��L�\Nt(Ԃ9"�o�t��Y3�;��w���j������`�E���e��4�e4^j��g�+����*���WB��cR���̥�*x*���S @!��i&���쏈H�:�җ����qK�h#'������\���-�K�4���QhJ4����@���D��zX���3��Q)��qv�Ta�1�n�L!'D0�3(�in/|�#}fzw��F6�|�ސcK�,��?���p(��$-���PH��"-�
�b~�;�^5�.�}��xJѺW�o+�k>ǭ+m�a����`���n���Qc9�bw8�f� �wNhԒ��y��a\V�J�2)��OKS�7rC�����P�بD6�; �:�tMg�����]=�IɏnZ.w�rSҊ*��!��M@'<wc� ��HRY�X���1G}��/�bL6xROG���,���R�7?e!��k�
�cDt'NR|bA,{J�����?����uB�+����I'�(DQ"�[#f�}XOo������a:�.=����uz���r�'ʆ8�����*M��<Qu]M%^6��LOg?�Ѳ�\�T��(�}=�	��zH��h_O���+�9�n32�t�ՏW�'�Ld;��\:Z`��H��$�g��Wmi��2���l��W�j�;D5g����F�I  �YlP\�7��>����+0�N�s��aX�q/��Rb�{�o�(|���j>ִ�>$�,�?E!(�!�2:t����8w{��9�Ё+"��j�ց��"�x�cŁ,X�D
F���?�y�X��w���T$sKU�{Tݛ]n�K�۬?�٣�k�:!�M;"�)���?,utN��Z����|��p�T]j垟��������G�Ȩ蠁}.�7*��Pt=�����8��.H�,k��࢈�ih�ŲJ�Q�wov�0A�� ��O�xj�ވe@k�w*ѸM�@��T��}O���/��0xddS���ђ�5і��5y+��?0sb���l��X��r�5徼�]���@씃f��j�4�HDrmX�m���5�	�U-3Լ`�yo�`byu�ݷ�����\.��6��.����LQ'Oܖe��
�M�.i\�7:5K4<	�&��n�$��l��P�F�t��?v',9W�I������00J��<ӳ��:�G;.d7R�\Z0]�2�E,��Dڕ�,���d����LV"��ho�؈��H��!%SU���z߆�/�,���=��i'0��S�"�l�qӱ.��DDS�w�5��D媎&Ee�� ����
�h�=1���箜�5	�(ڠ����8#z
`��Pa��C����6i�+���UO��S�am�L��Lu��.��`������GI��}��Bht0nۓ��;U�׉����
�.l'�Ln( �l�1ڏ��T�i���Xf��@�y��"-}�j�Nc�$"vgz�,�ǭ�
�QP�̭̜o��:���bq�����욈���U�(�iW|,%���z���a��T@U�o��*/��1�9�b��f�fW@�����=6<�(�r�a2�/d���l\Q�v>
�G�K���Y0ע$�We��kq�mY�H�O��F����Jj�gU�w�]v�p���p����L�/�K�m�����+Е���nE*�*��S�l��P���e���GFiW�")2�GX�hZ�Q����mv���;5=s����:R*L�O)��_E�)3���f4&�EVK��q�\�)9�KFP��S�;J�t(s���A�p��}�-.S%<�g��U<���8\�Y�ލ���r]g���R�Կxz���Ho�v�ש�·��|����FoE3_���@c�XH)���D��0�F�r9O���֠m��B$s���<��~���W�Q���!�%�Q�E�j��H�]�g�#�)]R�&�d�7�Q�%�u"F���;�I@�+
z���Y�;���7�v[T����I1r�C�vp��y'��(�jv�n�>p��,��g���`���ilFk�������4�a�T���k�lޮ|����	x6��sA�B�xs+�i�S?��/.�/�p�@�q�)"���+�.�̠V _�Uj����V��n�r���I�򳥛F@�*
���v������a%r�q��}�G��OJ�z� �w����c��x~HȐ��4��`����L��\�^ſ�Wm{��R�.�k�Y�2��zqkRԺ#��	��^/�!��g���Y�o#�� a�7[��I)�3|��fQY�Iz�7��������Zc�m�����w�T�g�cm-���Z&h0K�=��v�hՌ�~�uQK5I3R�M-Wr�pn�{�6&��h����>�0�7��=����W`�(�0���瘽�p�՟��`%og�M�~��]��s-H�=�Xw- ��x72_��K�p��[b�GY�i�{W>'�Ht�9+7�v⹈���o�(CE\��~�ŋ����.�/�d��S,Oq4���۳E��v��x�m�F%�8�č��S�Ŷ�������tŊ�D�[f�Ĵ���<�ц���c3q�~Jꖨ�L����t�9��Y�b}t�^�S��D���<�I� ��o��__1|��gehJO�#"�2X�O�G���7¤�0V�p���ұ�D
L�IoTRHxS�n���`�RR�GB��b\����_b5ʬ��C�msޒ�7�I���C�(Q>��\���xc�b������Z�'�$08�Bj')��|T8"8�tڕ���$J�}ά�Bl'*�g5����R7v��g��!n��]��+���A���O��Q�o;!�i������ ^�zRz[g�>Wظ��@O��wj�!����b:8=o�
�p�aW~87fq�1�=�J�?�?^rh׃,YX���)gV��0��}��N��_*�e�3�(X&B��D��x] �9U�:"���k�ʻ�ۻY$�A�!��:���I��V_B�|���.ݨb,��EXg�/(0O�u:&��@�Z��n,M_���ZC����Nb���#�A�S;.%�:G\���g�*<�������c,�ͪl����o3��a�3I{c�Tx���1Q�q��Qk�ݵ���%�U���T�����"��
�Vn�?�W?%~����X�l_�l��/�jA������u�oi��rr�K�'��L�{aX�L,�z	�q���e�&�r&V�SUIv��/X��<H{�����	w���/����]���?A��E3a�Ɇ$nK�D�l�5=-A�J�NE���,�M4���b��ė��w���'�y��M���I*�v���� tj
��u�m�e������f����.� -{!瓠*�Ұ*���SX��a�XSa��B�����}�}��n��<1'i�� ��nV��'t��$-U�Ed��S�l��W�6&�R�+���+6��8����E��i�z���ԲQ��o���\�wC|V��C�S����w�,@H�NP�)���lq\�Z��L1@0\�&���ˠ�_�p.���) (�L^���[�E[.�Ţ�R���1D��=�pZn��"z\�gs�ƍD�"*=�=Mڮ���.�u�J��ZK�v�Li�Tب��KyP���xe�h1NvpG�!ѯi�e�8	{r��c�L���t�	f��[�'���-��j�"�xݾ�6I��q�l��}�?�.d��	��"�皫�I)~�mj�g�Ҥ�m�`;�?�W��^��Qh��ǭ�"Y�],���i���C�h&�عqi`�*L�� ��N�g�t�I�X����fʔم*V�M0�h|U8-1 �9\n�y�˄c��%wˑ�|S`f��|�,�d����Fh�[�ǻ�r,>�ސ�5��8�VǼ��xd���/��|�]h��SE5�p��k,��J�S���J^PÕy"C���\�=�9��S�.Fa5䳤M�#���S75����۫��K�0��=��m)���֩����l3-1�*/J�u���?w��a��xXf&)OV�8"��:����W�SE�ë�/��7d�i�L=\0X����F�*Wp�������>�4�Б ��������_��|n��0��/�� M��o�B�ȣm:��ʖ���v��l6w���L2c��ܺ�1M��?���(w�:�P������2����߳���Po��i�ɏ�̞�_p1)���T�-
u����5Z���3O�P���顚��z��i�.4��1R������cY��1��b�[P����p�86y8G1h���ӈ�4B�].����P��몓Q�E:w���6lx"���7���?T��ڭ�t��� d���m��o∜���s$_�T�T�@gMI��"�����`^��iPx@�L�}�oIʺ����C���o@C9�i��o�'[�����v�lc�I?{U���o�SXS����L�ۺ
M��l�//��c.�~��g�$B2Q��+4����i*
���U�!�+�7�z�|\Y�h�y����_+_J\�p�O+�4��z���e��k��=��*�����y�_O+��⫞I����.�S�������U΋��y�G7���VG�qn}�ױ�l����a��W�l��:��	��֧�~\��@�:-�3E�э.k�F�����H7e�X�z3r��n����CxJ{��I���-z=a�*������*+���w����"IM&�y���j���t�.k�r�ushĘ�K�"��A�5%`���u���ga��84����a�z	K4���}`�r\�X!z`���*8VjY��[)��"�c����	�$e����n� ����������E�MP��s��U)��;S�a�Vo���F�k^1���ғ����N��_?��ͪ��/��[	����?ci�����R��mA�'�0��Sn��2��h�5LE�!���e���&� �M��b�t�~CMf^��Xk��Z��r%*�FW"�mJ��`f���z1~d�9��5ζ�*4(3��IHN/+�����Ȓ���fƞ�̋)b0��������4+U#�
�Q9�EܚcV��^sϦ9Z�1Pw�w����0Qx������J��-.i��$� v�E��i�5��W�)���ǔ�������訆�G�D�&���*
jNfÛ��Fi@�M�1��M3�-��3rk��\c�W-��@i�ę���<E�<F����֑D���c��>�w`_"�`�
X��4A��Frk�@1�a��mHZZ@��g��.�ye�>�hѡ������]>�`�S��@���ю6<"!���G�̈M<�C��!Ì6�rm<渜|�D�)�Y��:�o�4C�� � &
�r�������/I~ǎ�a�PU_���F�]�wпK'�<<ƹe��P:⳯͔�,^��:��>3:���|:���:/چ��O�X�$Bpg����hR����-$��k��7e4�-�"}��}iB�y��hjK���l2q��Z�'�W��'
��+YSM!�C�P���v�Rp�l,p�h�<����g�"��BN=tv�u2
6�5��R�=3��Gv�5o�L^^�hu�.({�4�+D1
:]���{Ve�V���֥��k���W〪C[���5�|��N�-^��][�g�_�c?��P=�Լ�CV�0�* y��$O�iŮ���/+�ꝋ )�'{&p:�� $J:�f�IW6���:��6��A_��ٴ��{c>��A��Ԯ����`ok߈0J�~M�߰��{Z�����P��E�^2p�uO���P2��R�l����;1����C֦,/f���+���T�v��8�[�8<��.KeuAj���ܼ-����--�@폅�ӎ�f�����c��G���C��|�Oi�����k݀:g����ʚ�/1'�2��\{h<��u��`/�JZ��)=��0���Th��
�8<�n�B0aK��S�Z>��^L�ΐ���� E��-�Kv]�������5h�,({��F7!q#v�@
�AzB�����>�DU��np�U�%��-)�d`P���X�}���T��\�V�@lF���^:�
�k��y=�?W�x�� �)f)mz  6V�
���6�h"����+��4�ڨ�ΓP>��`����5�n
�\��e��hS�ƴ�kl�.�.����s)\���#�hp�9����=���7t�����6���5����\D��$;̜�[8R9@���\�zD�qo��j�az�}��B�cU����tS:��u_�i���խ���)e������-Y��V瞺�!�u��~��ʅ�2,�<"Ic,�[�@���+U��	��0���ޡ�O8��MH(��6��Tg����w�3^MBԻ&Is��n�)&������ȖT��{��(b�������?%�[c[A�`�:pS��S�5���N׉�Gn�UE�G;��Qm z�S!�
$�����K�υ.k;�_ݫ�'���u`�������~r�Bw'��v��b�[s���@U�t�1��h�蒮Lmb�H�;�b�2��:ˏ�"@��%�����?�$��v�"���_��iT�c��ι�KY��	,�9��}��@P b<O�N���B�-:.�ϛ���\����Q��-�L�{��n�{��I� *��9|g��d�-]}?f~�5!j��%Z��!���)s�M�B�=X�Q��ۻfb(��f��,�k���s <|Z`n����*G�0��}嶼+DJ������Z�^�6���ZL��3�pm��r4�,%j�����J0[ҵ'/#z��Lٚ����H]:@�ӨB��=q�Þ��Q��C���q`�AHL������,����{|��ʴ5kW@�&d9�Y>^F�c�3�9����E�4'a0O��W^ND���I0��hD%��~.����1zqq���T�wg7xD��<wؽQ!8���Ţ�i��)��-^e� ~V���ӡ[m�B�,�m�8^?�jB�h��(�g�f-���=#��8�p0Z,���e�>�  ���W��Zg8�JoZ܇�\�-֡�KL��
��y�h�o���~�3R	hS�z,�����X��:y�/</vMS*���Ud��`'��,��@�)��3[n���痻��

>��{�9B�;�(��]:7�� ���bW���Cg_7��N��:.�t�JGO�^ 5�W��k��E���*�o�!1[��T���+Hm�� �!I�-]=�����nBq�e 7Ͷ�2GҬ�'@�<<,�X������SA���q>���o�.Km��:#9I�%{9o�^�lGq�LR�q� �M����H��r�; h|��
Z�'���M.��1�gT�D:�X�'��IR�z��)��}E�=���;�W��
�_ "�'FΡ��F$��_�k��MoˬLr���6�������܌2�dorYۇL!*
�-o���V-Ϙ
v���V��́�o�ѭ�ȧ�t@4L��J�$:�qv�=';L0���KZ���w��VXvl��}7���SpZ��8�B�����T�d)l:e���U�Д�+�n��W"�!�n�FO8�]���T �OTwE�ED��/�����o��"g9���y�G�_大�4����!�v$�2��R�u6���_��|�踻���.*��3�m蜹#y�������;3{�hd �m��|#�%'��+�<����NR)~/���Y�D
6���pw��,ϻ�x෷ش�^C�y�!4�i��]FQ�flѷ�nu����;S�`�b��J�];y�p�N��w�_q�#��v��}H���p�owST!JG���ބ�RUp9�o)��a�-��0\�W����焞x���yc����b�ퟻ����N9�2,{B��9�!M�bX��f{�-��$��1~�4A�r�S).龁܎��EJG ��Ub�Y&��?ĳ=�C�2/p��ub����q�΀���R���X���ӽ;k�-�O��cN;	��4z��K�Y��M�f����/bjE�γ2>4i7��c������]*����Z�-�rA�V���ײLJ�~m�?�r`z,��Cz��d��l����֯�?�s\�!^��j!�%��,�<�P7%�����S���H�����'���X0N�\�Js*� ��N�0���zT,Q����b�!Љ~z�B�*��1$��Z�سr�4r�D�w����m�p�Ƽ�~N�N��+�7_��eg�d�L��� |��y~�����5���ڭ@�F��h��>����ԉͪVV���#D�
E��Ֆ�H}>�M��w�u/R��uO+��]:�ؽ�^�ð$@y��������?��z}�B��8��>(�Go�N��iF7�k�.n�V;<��Q�PJ�	�9�k�9ĿK���N<��͕�u^�v��:dQIF3�K0Q!,�e��>�T]��T�:F>��-����*|�:{nj��#g�pޓ[���$pbM�a�?� Nŗ��.XT���t�{+y�?��S*�47����L��n���3IXl�'���RvI/�J*2d�p�mz�,tMR�����^�!e�.UjH�P��l-�F��?C����p%�=�s��pk����]��p/%�4����i!EET�ҐgQ�:�x�: �ܨ�=R�
��A�Hr�|��Ӑ�Y�󈫟�,�x����3�A��xzE;M�ҵ���x���5줥�o���R�闷���`�R��͇�����0�N�"���K�*�Gb+_%rt߅�Ѵ�T�,��`˵�B�|u!��H���,��Rq�]L������'F;@L��^dZ�`�b�r��J�|g:�Y<]K�� �;7��[�P�U`����D0��Y��;�)�Lϋ�M�g�ma��,Zra�8`+���yG����*.�(�#�$�1�c�{�c���]�@z�r�L���I��l�"��ǽ��lUے 5^Y,�z�C�/'�@3�&��&^�����ӌW����!��),�Μ��d/v��vڕ��T���ȶ�	��I�Y+3���\I��3Cp������xamf>�I4�&��X?D5���2��6��<) D��K�GE��s8�?�׆���Hd{�������抴y�&5�8�����]�7p�gA��������C�CY;>�Tu�������"-�ܝg�8�0�\L�*��X�(~$�������ץ�Q�f��s��̲[�>�iB�8ұI�gϨ�G�O;0�,w�{�59w��oᒧ��Ք?)KMc�(���+Kx� dq}eW���`��Q��Ư�fw�_��.�����b=$��}t�'JC���EU4+i
lk�9G/S�����Pj��3P�VU7��IOrt��OK6�\�EP26��T[U�H��S�)�)H"�<�@���.Y�XDǮ0��yh�UY�n�����z��R��B+�_�ʻ�E�C^U�� ��,9��/��,]���a!R�jT%��")t��\�ׄr�$e��Ϸ�����1ݿ�W>�$n�`cmAN�FWlيO��(��ǜV"��Խ��61P���\K�Yq�m�����nI���#��Ĭ&�&�õ�������$���ƽu��t_�8��N�Pf��ۙ���W_?�z��y���$wY�C��fp����kMP�}�������u�Z[��v�6���k���Bt_{�3c�%ϓOё�<�6Z �QM(��=��[?��_��'x|FMK�[���W�)�o�MUz^������9�)�rڵBA.��LY�}Łeܞ��߮΃!�N�Ď��$ M*����;��d�})_�W�_�lef����4	�6����Jm*ץ��
A���&�r,O���d�ĸ��~�I�A�S�Ѭ�����+�3ځ�����d�!o,}�H��+���,�F��0�/k�XgՉW�y[�m���=	"m¸*iI���DN�M�ú����xMV�%M�xͤR�)xN���%�n���v���+Ё+P^��'`F��-�0�����
P*��~��K��x�-���c�e�y���LOD��rѸ��	&9US�43M�[����B�y�L���v�:(k�F)G%Z�:�Kj@�����*޸r�eO\:b	��K%W�a�;�]ѓ|7�w)ҞfD"CC@?1���/���H�`f�ń��+r��7���S����^&��o��z�������>�  [�k��襓c/���28CqSl#B���8�2�� 1y`�P	`���(j��n%����I�f ng.��wn�lY:F��D��ͯ�����"\�wY���������$��+0���vH^f$�1bu=�(-���)x��Ow��ߧ���Ј����KܵP�7`�U\rH�<�W'O��zV&��ݖ7�0�
�̻��,?JeA�u���j�N�%2�| <�=�\�@-�
�����n��N���ܭ
z�LVZ��U�cc�%�v���)�`՟?k�$Z�H��E�<k���îk�jnX8w��g4�ة�~�����HGWaU��<Y�٢a��8�y�o�%?����{S��-΄ 6�H��3��KTbhG�A�g�B)y~B�	�">�j�06? $Rk)0����Bu+�mG~v}��П�(�o�4M������eQ���-�`�����Z��3F��v�T� <��[h�@� �n��YI��)5l�Ek��Emđ:�`��Ģ�+y�F"<L}=��諊���x�(��fP
pc�ʖ��&��n��p贏��F��~2�Xk?J�03�
��䰧]j���)ݽZ��j�� +E⫦ք������j^���WA��!�X���"4nclK�'T��wŲ@q�B�>��Gq=%�O�:���z>�Oʙ�0M�������;���I�4?���Δ�r�P���]y�/�e�ۅ0���VH�E��'~�F������b.��sP���O��!�OH����� d�4��[N��/f/�?̜o�vi�i��Z���P�t���7Ƽ0��J���6\�d���]�M���J��r�<A�+UtP@*�#:u�gz�ւ֠���VA��lg�S���p���C��[�� ���1�k��c)	�k}�2Q�VCB�mZ?J��5u�ޠs���)�u-pߔ�qE�´�m�q)WԹ��#Ќ��B_C�:���Gt�!��JRT��g�j�H7��O e�����ºl{aԚq���;=�O�u1�	$�D����`��4�Rq��&njF�߷j۔&�ݧz��F�ˁA/�>^�6��_18D�vP���PW�j����]�K���4[L*�ƒ�Ձ&����cU�����YU����@�/7�4�;�$�gy��e;s/����x���@���P0Z��\9�5a8�JE� 7���ДL���qx%8S`�L�B�{���4�Z6����7`i>=�ک.�C��r��Zzv�k�A�h��c��Ĥ��[�Z4g(/H1�����3va,2�i�����/�/�.��9����u�V��[TEĖy�m�]8])p�bc%��t��{J
?�1<	�FCc�0�h�Q�'q��AP�n����Ԕ���3%�Y&����)h��0�mg�m��N3��er��y<�1+Z"fׯ�4'&����r���2F/���e�k��^�"=����gO	�es1;�S\����fYZ�3�X#/�pi��'<Y��FC�H���K}����-�O����O$(D�C^!���+@�h8.��ܵ���x+d�����n.����ű@&� y��x���Ҍu_�ۥ�-��~��#2�$�P���i���!�D)���S��Y��K �N5[!�L'��@�	�\�z�{��c@�'�R@����V�q�D�V;�h�,�$��G��l6���>t����FU��X,2&�k�7����έ�������ǔ��nȓ6��p��!�My�����p�Cm�� �x7Tw���*+w!��'pTaC����*��_��1��A�ڃp{Q��=P>�k@>��W��y�<X8Y�f֫RL
xy力�y�˘��G�ӀS#:V�J�XMR�)�{���	=2P�����{�W�����%�IcK�(����a���/py��� �2��Q��l�}���M��~@[E��jG��1������*ȓ�7v���(,�
'2v�STSʏ�Y�v�e~u�?�����Ұj��귧MCu��ᣱ_�/��?e���ς�pЊ>y��Z7��=s|W9��7��)�re�ڟZ��K�Pᩆ��/iZ�%��� �rc�2ib/G��k=���|�&$"<*�f8�Pu��w����U��B���a#㐄 �?�'�V�[�x�$.��xTmX���y�ЭW]�ܙ�5��v�<`B(u�q�z�`>c��~�Z)����z�k���q^ >J��&�A
H��k�:R�%�@�\u;�n�����!���}o6D\����s�K+Gs�%��ȳ񫴌�н�o9�f�ݕOY���O^X
;���]�Z�M]|)9~��@���Kj����4�[�"h���y����m�A_c���H�1���7�[a��.6��;��	#FQ&1�Z�Y����.��c��S-�e����;p ��Kh�ڝ�OJI�9[n?��	����K;,!qb�:�$�k�ri|��v��^ָ�k��l�������7����r�5��|�����zO���i�9^%:�����>C�K�[��&!섥2�i�����)V{������V?!��v��� �^�*�-��+�t���6��]l�.}�y��at�k��Jz�.#��/K@���Szp�x�J6�Vd�`��k���=�/����8 ��:�~�O@��NZt�dq��Jǽ���"�펝-X�*�4D�C0է�}�K����_3�<9�\E(J)h�jҐQ����9k�v��a=��]W�2���殮F�@��U��+�R� Ҿ�v����n,�'T�֩2��=� ��o��������~�-$}4���b��
Y��w�E�m!�iF�D�����	�c5B�|$P�	TX����k�gW��.A£\�*��J/Pݳ�����{|�9�z&J4�qj�i@� *Ҁ�P������1j�:IlO&�D9y�Wd�Ltޭ���L@��#�a)�v��W����OR�# 1 �H~���f�\s�m��������e#��(˛��D(����}21%�b����j�����H��#օO�bm檩%�"E�W��jG�i��Z'eB�s2�~v:��h m#�W�y���Y�U?�����ʹx[����1A�Sׅ'2�G�^9k��GH[� 3D��(��3P�	^"�0�d������+$A�H�5�U�Z�*h�>�
w�J=�a��`�ͼ
��&0�w(�'�N�s����+����do�����2�[7���#u3����>� D�甋M-�]D�=�:+�4'x�䝵޻�H��r��o]�c �_i�����ܱ�/0�:�@+9b� &n] �߃�F�G^�&i[�~��ھ�V�%�
�YPWܱg���+�ب��(��9t��j�%�b��g�4x���g��U�8��P�ϫr�9�������j����'���qu���p�Y����-=��W�ɛ���U�?��	�$F�7Vb�}���V���/����(S.̒b����k�����+4�=д-�~B�c� s�V*��r��z/��"�:������Pa��ّw�����IW�
���g��>��۵��Hђ��x�v-^�H�����ا������y\�k�U��� �sd%�d�_�>_���E��mB};0�� �����g�QT�|A���5\�uΥ�s�^�X���gC���/\����Q���[�/}�b�3��z�[�/��w�ڕ$��4��o�����W���'�eL�z�.�������Ӽ��7��ded��5CZ�$�W�ܧ�� �����:�G���E΀R�YEVg{^Z��E;E�>��l@��4�v��,hS�o5�+PeUW��-�N<l(���΢.j�jq����ZrO%˖�5��.�=|*0d��^(a�J�t�)���Z�dBt0���\S��|޹h�?3]�IHb̲����~wG�� =�& �)�Pm�z�������)#�5�Ǥ�ԭ��Fa���E�s�]�O|G���B������>�
`����&�B��!b��W}"����Y�R���9B��CW�Q��m�"{�A �h���&����.qeg��&5N���r�<��6���5(Х*ڰSl�4U�����#`���5�zۛ�ܒ��|3��� �M��M�k{
vB�X]���
5�y:��Hy�a��_6�/d`��a�!Xݟ�l'_0�����E��|��!X���ͥ���w ����Dř�r�߆�Ɩ�+������Y:�JAY=}B�d:�$��T�$�'@���z����e_3`� �u9�F95���ȳ,X���-c��b>5����2��f �u/�o��c��(G�H'�f@����_ ~�a�`��9(��>$-�K�k�j���a�5��PȢe��b��Fޓv��L���(ُ�����rLg���S;�p��,".'0<�����%E�p,��&	�w)�jb�J�Q����=��=����f�|����ߟ,�bt��Ö��E��������[�n`ژ�H5:Rj>�6.�Ci��/�\�m j1�
{��Qp��q��Z���l+�^S�ª{�H�p�Q����������"�ǈ�qp���X�(mF�M�#i����W����~$;o�-ġWĭM~���7)M7 O>��u<��W�e���t��5��] ��O��R�C����`���]���	JHn�*qjsyr~�	'4	f��<3!�[��8M���F Gύ1<���a����������t�Q�cɝ���z+����%_	��3�]N.9��_٣H����Zf%��!\�H��NL@�~�w��G�,̍U�kL�o�������p�+��F���j�Hz�U-"��޼���b�C��ml��K�5���\�帢ax����oZ�ۯ���$�o�a��k+���5�!��S�F�4�#���8�2���f�!P
�#���iV�Z��#t� t�Џ���>.�`GYMQu��U�ٺ�ǖ�Τs�}����P��`����DR��L<� ]@X���^�9g�"���B< ���nT��R]6�@�"|�b��
Z�xM�?r��yx��U��x,�C��6�L��}#S4�����N�u&�5Ñ�`K�.�z��i]�0$b�i)�>,x�i���❁�Wn���8��c��V�c����+�A��oѦi�1 *��J$O
*F�+������닣��xR�q1���A��g�N��`��9_��`a�3n�\A��F�1J��b��(�<T_�Z0kXƜ^q�e�+�x>Ek���9��v;)1Yh!�ҿ<�{��u���_�D�������s_�;�����҃D�1�7�kR�{V�OB�b�Ak��8��n��Z�Ύ�Q�fcg��ɰ ����,4FA�"�a����.L�
��dD�-:c6^7N<�~�L���F�b��U'����M��j.K��Npz|^�8Xxu$��Z���u�FN@�F�Y���^���O�p��^� �Ѯ'��)is��*��$T��o}ȩ�4/5���:��!��^�%�*���PQ��󸉊궷O�&E���}�Le�h>[����_�*��c��[C�0p�2�/��帐�I{�i���-sZ�[��V��-E�L;�&�
�ߊ����O���,�鵡�(h�:��
U�.�W�����&D�d�Z}ѻ����Y���z6����W�:D(
5�W��8ʶ�@�襏�ET����*8=��쪴q��^�
���x��%>��xQ<P� T�NC;"b/J��ݞ����Y���_2��D��L��J��~ͩ�EUl]K{�a���D��vFA~�S1�=���,�.JQ�hþ���ݟ�W�����3i�J�WZ��k�!H��;��ha�D���wֻ��t����v6��a��ׂ2����%��mM$&3����Gvx�H:������[uT;���Ug���1�&�.�}�uQOrK�#�-'�%�/M�@i��z�9�U
uhG�&:8K��_���������.����ަ^�ke��fp|�3[�q�by��/����fۜ�4����ݕ_ddv��������ARW܈�s؈���.�Q~�y�����n(���뒸{�.�>���3g�� ����ނ)��8+��l�
���ҋG��'?o�;n���.�=��Z	�H�3�����w����>�#�9�9���x���7�H�:卬^k�_Yz���(�;���1^9������F�/��%W�?Q�*���$�bu!��{޼�d��ȭ���������	|���J�"�q?� �#\xo$�ď�ܖȈÃ��:��^W_и`��6�V�����3q4��A`7���D��Vu5w�y���#F�����	<� �Y݀?��AN|���ӷT�4�㛗U�`���0���R>�ߔNs�N���0b+�Z����˯�	�5v�)��z`�e�	R����x��e�^���a��~F����ĤE-�L2;H�3l2�H�?k��~<i$�-Z��Տ���!ѩ�H���n|�F�C@Y�!���j�@�%*�7�#;���N��Wd7�iHg�ϟ��@Q�N�-o��sS^d�WZr5Q�!��$�+�S 4b2s��tw#|��Ԋh2�{����M�fӦ���~�Mz�	���}�0:�Bi�5��H��|��Sr�w������l�:��t�q����9)��
���T����@<�;Z����n���w�#hi'{������<iŐ��d��c��/y��g�Ȩ��R����I1��������zl'B�P����VP3y��r̢�v^]�~أ�N8��p������&���3�B/iq�]��ٿ���3頻&��}?r�Cx_������E���%���ğa�&]i2a_�4\�0�����D=E�6l���u:3��vQ'��p�EJ�����JH�����vp�X�Qúڃ��3��bb_��]�h�5?x��x\��p '�Jч7�f3�+!pjU�'6�s���_dk�~{����u�u����3�E�@�!Z/�u�б�S.�8$�j�d��R����h���TɅ��K�#P��,N1Qn}��ԋqQ��Z�&z�99Y��)hc�D�lo�e�$|�5���?��j���+Y������Ϛ/��T�֥�h��n̮g��.��<��5S��>��9�y���<WrpZ������ΚA� ���j���ᝉ�1?Ma]��S���L|�%
58�恃x׷��M��ˇ9���g&�L�>~�W��x���V=�_ ��׉9'[�(�ֹ	3�ٚI��5l�?��!�'�)���K�yUZ_�`��%�1��8#v}f��2�����)��@_0!��q��e	�u����hK�Lh�"i�/�vb>��;FZ$ g�O�_,��G:�˭-��v�P5�~�L(m1i�$ϖ�v���b�2��]p���?��a�)��m�(�L������Yao�#ΙH$X('�僕����� ��[[\̜��ok�eR3g$�qV߫�O��`q��3l�߳W��l3tk><D�|)�7m���%|��CA����js\ؙ��)������J�������PV� ����$d@9kF'\��b%�t�N����?�F��
K:9c&�ٵy�^˟#�'z����w����k�<OsZ�&�r>�F[4�z���h����{��:J6y]���$_�<ĉٯ�Ij?�����8�膰R��
��K�n�^j���RV�I�sW~1���*�q1��1b��3KG�Hu-��߹�R�,5D�v�����93\[�Ui돀S�7ֵ^ݖ���6����ӎ��%�'�#�����Zq��������}�.]
j9K���"��*����&q�~����g������W�Z��^�~�
�j��T��aRsj�Y�7�A����Ddi�|m�3�S.�`�2���������I6�说��
�4J¢���-�A��,��ke�Kpz�Q��n�̊_<�X��G��sF���L���]8�t)��ڗhT\��՝��h�hS+>�0�G��3���`a���Pɳ-�N_��������Xn�n<$���Ɗf����?����b*J�.�>ݽ��趚�]�������J�BM�̄�d�&���rհ�͸I�����p<���T1>��<��cH��)�O�1��#�U�b��.-�OR���L�Èбw��,<��r��(��?� ����d��^�W4|��ū�c�!*��j�%���}�Z���+m�Ho�$�qU R�W*��`�o3;�+ذa��k{r@�uJ7���2����bF*��j�ʈ(/����ц�>B'�O���"�ǫqtQWC� �V`8h=��D�p=t9%���(�mYE���>�=�6��s�����s�~�ρ����[�	ea!" O{��'��F�g��ށnNx���x�O)���U���ɜ��ڲ��%���6����S�I��y��4�jV�DP��q|�j��� pd�(@�zw��u!#���V�֙#������W����4��t�w4S�q�{���.���,t����f~����8�O؄��'o�`�/��_�C�xB��,����n>�4xz >�/�~Uj��ЁÜ�l��w$SZ;"���b����C`�#PY%�4{�����������%����3l��|��'�Îv��C\F�i�a�|�^���ɣ�e�J�?Q������c�<�*�9�
��Y���,g�#6\w4�iS�}BL�n��+�۫͞L���Xn��}���_y���y|�3!FY���F���7� �(��̴��EݲRA��R7eQ�Q�y)ެ�4�CRQ�E��v�@U�8g��Ⱥ.��Bz}1�iA6��z��:���BP���'�z�'��6_��[��k�b�2���'ŋ7-�vƀ�|"n"ӄ[�2q_���vzy]��}E��@@/����,N>��z� �58g,��D<:�`X��x�H#��ן��+Xս�	�U@�*>�Q�tS�<���	{�쿑��*d�k������0����D�^Y�{*Q�>�W!�E7�L��x���[��>Ad���Z%�fE	K�7֎�`+�,[<�h�P!��<CkL6P/�:y�>��q�z{z_�%U���.����H����e��Yoc���Xa���S�����|�l�(Ѽ�A#լ�nWzm�C��'F��ݸK�j��V?։��ӵ ��}!�������)Bm? Cp7�8�\5�`d�mM�"��	� 
�����~�.�-�W/��Ե��F��z�����V2�6�'~=/�tK�3���}U2�nD�%꪿�aV��cx��ҽ�hG�LS����y�j� �7@���M��B]�e��)���8��%�ӌ�]`M]/w:�E�G���ž��[=��WF�,���Qf����m���İ��h�`���pOKޖ�:�[Ƥ�=G����ӕkH;�s��T���<wr8#���^�M�/�?d1�,=���r�w����	ޖRMk�s��=���w>���M�<� kP<Cz	"�e9p~X^�(����)R��A��an#��9k�p�gV���m��y+U�����\R����x�����^���ßFi��9ѫ`r�~u?���>fL��$���F�A��,����\d戤UH#}�ͩ7�/y��s8��$�U �k!�9�+Əgt�9��`?�E�28 �	�^p�b��N�����-:�94�3��A��j��K�&���FXA��������ؑ:b[�yn{�oy�z��-�#��I������A�&�����-c	x���~B^�O5���/I=$�N8��<Ҵ�6��1�0�q�:Xs���	}�C�)����[��ll��(~���^�^E��]�]�1G���a�h0�%L�X/^�<���F���f�)8+5û`}�����4���	E)X�=��@��?�5��HA�z2���mu"g{�Xv
 
>�y�ߣ��6�9�s�k�0��G�a�$��`uc�P����?dŨ1\�Zw�^��`��#�U>q�f��<;$5��ǧ:�|�m��UQР��>.�0�|��i�z�Y��$�^i���w�D�I�h�e�B�c7q*=�r�P��*!���7)���@�/��R�I3V���g�v���jr6'�U/�����5��H�O����{v�?Kx�+�d��BI��zr��Q%��M��ūK�4@���ϓ)���D�`hƖ����|�{Gg�b�Aߊ�/����E؟�x���=)-�Ф��&���k������8��V��:�E� ���m֙�g#Ӵ�H'_��_�/�b�O��Xf%%txA����[�j+�ant�H��ƍ���q7�g�l?�=���C�1�kCD9�N`����3�,F��* ��v�Hn���w�S����$f=V���r��Q�C�Ι�ۜ�3�c��V�s��l�.j�����ܡ�;��yV�U������~�I/�l� ��B�*���.�Yaz�Rt�bS�
�����'��l�?6%$zX�l����j�a�6q�r�m9 ��F���n҇�����s\ŭ�f.����õtln� �@h���EK����Ƙ�m@*��xPx�~�g���{ߡ��6*��Bi*EIF���� �nhS���ZaH���K�tv{IUFK�.[4���낞�W�`k�����6�6�p�Jw<����*��}������-���Io4ʶf��!C2}K�Ԑ�Н����(�0{��ʨ�)��xʓ��
I��x]�v時��(�\dC�.|</:�W�q�8,���|&HlJP�-V�r0� �yf^
~��&���@ ��5����+68��;-�Zgcw�{�y`�����16�${��"5�f�[-��W�����G5
cNoR���S+�K5F�?��:��Oߤ��`V4ŏ��PF�J'?��)]����j�*jL*[j�|rn�;����Q�Gԋ�e�6�|m�uKR-}��1W�!�e"i�?���7 ������F<�"/ }i�)�L��rO9���;n�o�*�XaT��n����6
{;�fz1�� �N�:�4�h<	*�!CD:|U�:�
M�O[�]���[��ME�D��o7�0�#j�����^� �x�X�L�����k����E���[�r�s4���p;����8�c�iשr���}�鍬+�q���nS�y�G	w�V��jEV67�&S�X+[��}�~d���*.�	�8jAL�ñ#��ӑ5p�`�/�rC��m�"�f$��%M�
\��ݮ�}ߴ�gVQ,3g�^�$��G��	�O�r�@��,��R�s֍쉗��sC��ߐ���A���" /W��5���Icwvn��v7��.�|�g^��Y��#r~7d����xw�us�v��u��2�V�UY�W�#9��v�L�
�p�ۏ'Ȇ�=r@E|���M��խʤ��d��d��'�;-��\���ý�$�*�T����F�~�U�|T�mK�Q@s$����W���x[�nY$G���/��Li�kXG�`���c�%���=}���j����H�h�e5s�c�BsS{::v���*��ze��M�]�����mmO��Cf<9�f���2�����3ܢ|��)'uж��.�8r9�An�
�R�s� Y�;����4����V0�4�g-��ѣ�><�=��O����W�޳�9�xp���
�����O�^՞�1G���5�S�.���]S�����M�i; ��:�@�uۘ܁����y�'\l{p~�W4��ڍfhf7ն�@����.�\� P��B-8j�+��څ���6}ډ����N�Mss��%��-�`�Z�1���9�}ʐL��$��`d�
1g��ߺ�v� �K�U��H.�b�%�S��B�_3��f�ugt
v\&��d:���
����m=�	��:b��䯹79�+��t&ì���۱VW}����ܙ���Ӎf���-�Ǯ������G��-L�_
�sL~�߂T�;:�:h��YaK5�m��ß���;���d�w��ô�#�,̎GӱI��G�#%ơ�0ѡd�1`;q0��b�g�6yk�_�b����f!{g�
7��z7�MK,%��$�;)\.�Yg��9 ,D{�n�<x �e2�S���b��+r��*�̒w8<�����?�=�Ÿ��D,�93>3�+=)U�/�}H�EYaמ^A+͓�q2�`�۲]��8������:{���A����q��Z�E~�@nu��q�<�9.�^� ?؄!�o΍�&��d!*�3b�6�:6k�vh�8�!NG&bd�Sx��dz
��'S=T'2�l+- Ke�!F�0���Y���N����NΑps?Sw�35����Q��ث4����<���d��F��A&��=�q�ڧ]�pH����$Q�n��
e�y:{X}_2L�'*��o{���׿?/ᘦ�ܛ���g���,9�+O���!��}!��I\�ݚ�yH�c'�����J�E�n�ɨt6��O��ذvE`W$l5����h��&C�_S����(���xz�+�Y���7`�I�|~r�Q��v_4mc���ȥ��Dl�R��n���ϴ¡�N"��֞�ML���R��)i�����{�;Y���g�����ܽ���93��6�[r�+#�r�L���nf�2�ځ�o�v�T�a	{�P�$ī�g�T8No�ҍ��^��_JI�@��ǃ�m����슮�0Wb�G;x��:�,�鶀* *[�
!!݋T+� x��M۞?f��F�O�n��d��#sN��XG�+�:�>��m���RTR:�64 ��=e��M�3cʰd�t�B��>w�)��p�HUy������ĕ�J���Z�HA���3�/�ō}��Vp�D�Q�g�Z���{�-����E"�.�!eEvJ:�mKc���/�^}�����o��-�QM��20�f�%9����G�G�yЈ '����i7�����w�,J��<����M_���<r �x]��Z%�	���p.z�<��˥��z\'^+I}����>� ^��%�Ĺ��{W��E��7t$̅���h��<f��=��)���}8�1>g7��S8�`���ZX\�(�i+@z�,�k��z�'3Й]i*̊����x��!u~�B7�,�+=����]A�}���{���X:���ƪ�T�pL��.�u	(���B�߬W.Ow�i��]����+�R�n{��bḍѰ��㕚`Mꜘz�O �!�r��༳��-jӰXL|��P���nb�dc��F=�L�֙+!��X��D���������A������ �z��|<0
?��M�M�$�s����(Vӿ�IX�^�����/�D�x�緞���-c���B�W&|���g����5����A�/`Ӫ�}J�ӥ'@@��Z�$p���<�&UvIPr����OB4d�9���mV��|�)�^o��i
�cd�Wy!��?��`�V"�!��c��7f�ĂZV)�9I�/vo��7�,w7����9)F�_�"K$�T���a���f�_�Y�!�B�x����}e+�L}�TLk�V����,.�Z,S^:�����&ۗ�7��A�T+����T���Y�De���ф�<K1r�KB%et~���"K?�8�^�<x�zUN�QN�ő�?Ȟ�m�T�^K�V^�q`�%u�N���������v�lM�u�:����Η�Z���Ą�|;/�6	u��9� ��<15@j��t���]+1u��gZ��LZ�JaT\��
�(�D��QD�nݙ �ݏR�|^�@���G�UJ~�H��@��ņ�dZ��{�q��Z�W�D�O�1ci{��(>�wk��l��^�\Œ[:���г	*|�[�&�J���U�&\�k�4���8�֕��'��g>��B��Ȳl��~t�������ڎ=Gں!����qk4��vOd1�PW�K�6�[Z�V�H�h5$��x�F�T��@��<p�8Y��P񘺔�i��_�����/�0՛�x���jވ�[�Iۯz���Hڦ�T#���8T��,����(�t��O\�a���U��E�+۽��\t��/0�?2pC�V�4m �R���w ��6�Q9Q�_����>[]����T�	П��}��y��W\�rEų����`g��#�e�D��h�x��:�Zo�x�������;n�e.�έ�=9rI9���$޿Z�--���K�7��P7J$���J)�K���ن+57�!�1%�xO�a�w5mMx�oX2�=+H��$,bM/4ܥE����o��ߧ�
��c(�zM�n�hD�'�����w	P�����D����x���NI��q�S.��@�޵|�v$�4u=��i?�c�g�}r��$��(��U�3��<R�>E���l��;T��0n
K�&�1�y�/���>Bǂ4��r��bF(��U+f��Mj�~(5|��Y�e�>l�3"?sQ�E��U��~'W��3��U��	,�Á��=��j>tR���!#�}D�&�l/<L��O����kՌ;L�
��.�Ț&g�o�&=�9�g�ŧ�轙\��C'�3�$�
J>������Ƨ���g���N��3��e�z�M��#�\��Zo!m�2)?��{t��@ʭK�+0�~@G<�Qs��iPq��|k�T�O��q2���ʦzM��cƚ����T�`1a�氒�O7̓��B��yD
;NJ��U��Ó��m���ͯ����tk�U %��(i���s֋pn�kQ��W^|,�A-aB�E�3��a8X�����',�Ӛ	��蛬>t-$�&��K����Z��[!�F"��
���gL�S���j�i-؆��x�sl��<��	+�Fh��7���[�66�Ғ[	�:��������NŝG%�/ ��0S��}lGN��
GO����Q���cL!�F۰#��H+�r|�O0$�`*�n"�)��F5��㗚�;�/�l��T���k�ل�P:yP�'E��#�i@�z7�����j���m|7�a������/PD�ߺ�c��(U���J4��+�Q�?��ZL�\ѹ*r�����c=��$��=�Z��)��4E����
�\�T�4�<;ʜ^���o���~��̈́����`V�N�{˹�ӵ�f>iЋ�����^�����w�L�@�sν$��^H�]���֦��ܗ��������
��o�9|١�P��_e�j�$e�����9i3���C��W�a�"�zd��/C{�q�$3���j�֖�W�?�ՠLXl@O��m7K(����l�nP=�Ʊ޶-)�2h�"`��4���.�cn���DF� '2���x36� 5��0ך�@b���E=;��S����2CL�+p;x�Z�T�`v�8;�Hܔ֭4�3���p!l"!��	��pM���W��:l'#��v�+L5$��8e��a���]o���j��jH|/얕.�OU
���ywZ�8�l�:���'�\�" ���$tU�%l�o�g	q������v��L�՘�lX7��^��dܳ�:�CD�׿�g��n.�� ip�R4(��r��m��L�݉3-��x����_ǫNI���/��5.6�9�p�)��{!�&zs���wтs{�3cכ��pH2�v�N.�T@�K�%�aE��U�U܍"� gg{�NN�;ӆqz�0O|��`W�E�xHɄF$9��M��/��&6P��\{J��ϋ�
�H������������6����H��뱷��}���ʃ{���e`r��fZhZ{:)�t�ở�jA�{������}������J��I0���`؛�������8Z�Q/�>����Q���`�����	��޷\\|�-:)k���=�Α�My�_��*]�f��*.�i����c4|��sy�v��~�O7��P3�7^鞇�4�@����O�hg]9:g�a0j�H�E����-B�`�Kqlg�{��E(��*���A��O`�B^wҙ��t-*ZRhYf?�Yk��H5���4�:�Գ�"w�Dl���8dhq���^/�Z�Q��6��õ�2f��;�k$ME(�t���i.3b1
S^��.+�L�w�K �a��7j`+|� NV�8f��d���l�|�Dy�]ꕲ�v~���ʩ{`��ST��J�Q:�mG��kC��VIAk�������~+��A��'X� 5W�j���忬�ɖ�Tu�s\�aq�d�
��c]�P��-�-VX>-�܋��Ep[��1w�6A�P��E�;/�ˬ]Ow��p����勎A�	�[�U�������`�S��0Á4��l88ֻ���iPh���M�O�h/湇E�"�(#q�*^7��l�qnzy�)�B�}�A�4S �>p���{�R��6��5��w����-f
r%��i�Q��2\٦8&�f}��ui�����?�t�����yʋ�ۈ�	�����Z8�t����N��:n�r{��1��k*�+�"�Zf�}`����Oydf��(��?��qeJrC4�@m	ð�)�1��?�z��ya�we��#�����M,И�h*��R�ID%c],'s7��k|���p�,U��ªXCǶ�
1Y��3�a�ԕMa���xQ�<1�u��"�s���&���Ǝ	��#���M��Ȗ;�z:��Nv]�m�/�D�x�X���ˎ��BYWKy�Ծ�ZW1��#�C�8>N���kք�M�/~ˈ+?�8� 'vJwD�Ɍ�\��q�$�����L�A�+��2��4�h�^���eY�hG}��?H�K�ҕ�P�T�x���cK�-rO��a&��^�ojL+���]� �-s�a����9p���Sv{D�	������$^�mi�t��8�����W,��G�x��ޜ�� �es���4��~��Mq�zm�X�y��=G�7�!�e�Z#�$�oL2haN�A;��}5�ʿF�sl��N��ra6�o�wǓ'����L�AB��B8�A����5M.}U�M���#��/��>h� �.ANl��1�)�0�x����q��c�)vV�tY�y�	���Aݼ��&rB��J ���I ũ�� ���Z�[�ڸsd�g��c�[�Ռ>�_;�=E�9"|�!����"��rR �h�,����'mn�a�@G+������vɭW�qaw&��ഺ(x1"JR^�}kd4$�T;W�f�#�m��Z:��^� ��-k���"�����5�e���V�4�3��K�u��I��	x������vD���Nrة�?v�H�XzH�l�94��W���65�H�ߏ�Lf�Ԓ��Tܔ�ʝ�I�����4��c�l���E��za��s�1��`�yOǠޞ�����!�J�DJ(e�Z0��G�쯿2��RI�}>uk5�����?����,�r��g
�[+��E��p��V(w�Ӟ�D���D���I9�6���0��;Jŀ�:%�
�mk?H\�*T��ʨwL�/ ���?jê�&���I�c�C���Q/����	R�#��M���zQ�T��B �~,�/3RKT��Hv/��#cTp�d#S(�8[~Z]X9� R~0�P�2 y<��orK�>V3oeQ�L�5��HNVa�3�@�6����~���oʝr�a�ŉ/�18��eԼx�
1<�U��rBZ���;8V��|i��c�1��9>c�'���K�"ˍ���$!��!b�]b�����v��DX�&7��5q�e�DmmrYcb�q��V�m��c�L%��ǳ���?bқb�Ǵ�8Ș�6K�D�W��z҅�
Bccu���m�=�����3Y�gX\�<����5���Y< ���
+ ��+����y���;�]��ie
NT��=����b�_�O!/ѨX��n�R�k�����R�O,M���i��#sPk���͂�-T�`�ș�#n;u��̄�����*��h���B��#8����92�r��JطHO�p�a)g4+Yt.�Y>���������̧��¤A���6*�
T)���� <��'{O��8���d�昍�1옔�$�
�*�x��?�A/�S����$kh0���8A��
�"�8I)A�Ky�P5,�)�����z*�UOI� 5����م
�s}:f�@'�I?އ7�,��m?b�)�#=*]DI����\����j��`�͑x#��/���U,�u��U�-,q�����E�P�\�iZ�2j����)w+����x�ȱs&PX-a;l8��BI�5��m��>h�6vHA�%K�6��#��Ya���2n���G24�b[F�u���G����ʻ�X����v��,Y��zJ7.�B���+B��~�"�� �k_��
xAbq};��0e���I0ƞb��u��ǋW�Y������)]!7\�Uo���O��WM>,�W�4��������L5ጠN�Q���fAΌL�:U���>S��_/�*�'����{@��y��5+�G�Io�R?k�Ď@��No�����T�g��#+��R����b�=q�Pm��C�54�pV�z��s��E���MQ.��/��`O�ۍ���76l5����1�͸ߪ�：��=� �p��1*Pu# ߶���/1��OU¿�.�	?4���r�x�L�Rja� ���8
�D4��o_cs���0��Gz�q����T	�h�L��ߓ���@ygCM�7$��)�z�#��0�$����Zm5�7��gFxzݨ������R����Nt>�!���:�Wձ|\l��
|����V�pj�9��y������?�)1*T�î��Â?V�}H2tZs�M:���z�m��;v4�nF�4�Rn+�9������nr�Cv��DE
��	��j��&�+RY0p�1��i�vۙ�o��=���4S_��B\ ~i�`�\��x5�O���Pc
)��a������:U#��*^<�OE����<ɀ�2��l�w�by�Bn���kKqeX,1��M>/3�m��{�MZn���x. ����G�K�7�6�NC� �D0֌���������*��:7�5��r8�-�e@�)��M��Z��?������W���0*5�gN<�鶇��0��̓������v�!�V��z���K���i��Qo*<������FÍ1����O�>��r{�@��ht�����  �4�J��ݢ����81&·^�2���	H�E�s{�l�V�e�ݿL�j%��b�{z�L?����G��Z���\����>z�\�ϖRS0�ma�T�Wq�O<�a�z�#x�w�I��\Qj����˥��\�D�7� Kr����u�͢��ŏ܃t䩶�\3u1	_+�5����X�1Ym�W�z_��7&#�]/�P�jN#���s*�xu_.Ny�g����/`Dm�-�l�^�k��%n�ϰ�C\/�0�������)O���ν��l��r�_tXS�i����Y�R}ٟ���n��E��Y<M���}&�)����w��x�E��Py���I��3b�vT�oj5���>�d2�9��V�F$��)����U�E-��z��@x��S/��m09Em	�
��}m��ڄ%fް�&��O.��9�֩�C�8�o|X�ᓧl"� �ИE7/��G���yp�Hg_m��0j��( Y' �1}�v���
�g;���'���vq����c�K �?�ޖS��^�a	e��7Շ�������B�M �~��ۼh�G��q�P[\��ۛ�+5D��s_�����S��[Eh����K���{�3�sS�Vn�ް.���8q��1=�ы{c̶��'!�v	5^6n��o�'���B�"3�B���:�ࣹ��;�LaD��$��h[.��Prۣ�l����	��lDLG����A~ľ������>�Zj�	W#'���`1�'��D���P!��&�{�<O�a,�m����j�L���H-t�Xw�Ԧ`�#Z戵���c�cV{�e�Km�T��es��{9��C(S��?�቉��z+h�'�_��P_9�������3��-%�+�{�:��|c��O������@�j(�paUn�
)�$�-\�:��T�a�U���z$�sk�jhp����z8r��5��2d��5�+[-��J��/������ĮP�-��=S���Ms~����J�
R�*���t&;����S�w�Sq;ׄ��CZ�8i>?:��9�ȼw����?*��µJc_���
ÝI�L�����^���/���e�Ο9^���M)9:�:䐄�5�g�՗�Gٖ����;\���U��u�j�@l���DM�gs[��gɿ�5��j��vgY���]�}a�4@�wh;d�I�j��"��8�.\���%��=���h$�
U
A�D��O����#�@�ţo����CY�A�^`�
���j�B)�ۤ86��2�p��o E BX��4�����B�Me[W4��ZM�ʎٛ".ZbT�+?�g���lΈ��p�����;egrPۄ�����n֋5���ﺖ��N�� '9�WY��KЄ�P��xX"Ͱ��s�$1.��ڏ��!�fkj�=���n�N�8��)]GW�:�p9����8�2/�� `���=���y2'��A#���EH�\���CF���>9��"x�O}GIQ�A���s�vI:	�$ƀ�
 lXfG���Z��Lh���"`Mӝz��\!zC̀��+F�4�킨�C#Mq$��\]Ul��o#
U?<��`2����%����:�r,7�ȶ.��V�2��0�N5
K��h�,��"�XU�d����+����*!���b���i6Hq�/�فG.t�9��	vq6ܰ��07��nj��+K#�Bf=5�ޠzkׇ{4w����df���l�%x��
�'i9���l�b	��x�(W�T�.�O�{�P̦+NԤ�69��%��)@�2�4�u�R�_���)���cw����:#|P��V(����!^�@:W�D�z��MC�]�<#bvw�$�J艳Ey�vlf��6��2�5����Cϝ9�xB�#Mz̺'ڎ �E������.����6��<�Q�O vqD�i����U�*O?S�|_@O���;��S�l�N�X�~�(��a�a[e@ߵ���N��4���8��%ZuQ���<��\"�]ǂa�<HH�ΏT�mLR��<y"匩����>LA�񖕀� ���L��N��v�T�_��R���ݸgQSՎ�qIss�Xdx[8��I{F�&�����"�xǘ�����O�5�ޜ#2[!��0	>���g��y*�3�px�،R�`d�����l'�m��CE���c�n���DVI
¤��fM˯�DahuK��-+�6��=�ܼ�G�n��>i�f�MYC�p�r�D�����O�w��U����g	�w%����J"?��C'�]B<��a�_
��ꉦ4��A���6��l�{E�xҚ�+fƸ@U�ߡ��`�;1w9���!D@�,�P^�;��`?�/����Nﴇe���<�Գ���7����ޛ^ѕ����y�ړ�M0��q���U���o�zp�b+�����vqUF���x�Y�)��>@ngw�󍦮�&�g�"��Ց�L�W���J<����Hە�������oƞK�vq���c�������&T+Þ���s��=	u���<��KH�<�{��#�����lA�BSF�
w���܅��'L����c3�J{]�b/ol@B�R0�棽��%�G�[^��t��mՁ*((�#���a��ka���C����ņ�e*f����s�v=@aT�
�d:�jO�U�5&�O���vC䕀�˞v��QExx͏ؗ��r���5	��Q��`4���r`���J��Ud����W$sR�f��%6^�������� �f<�v����W>����V�й�\mK&�ȅW�����}O��g�=WnO����KY�C%����S�m*��*zՁv�����\�Z��,�^Ms�Z&6�ɴ+jH��{5z�X��_���0�:�f9�D��D�#q�3��W�D�X4`� G��pg����%�>�&d¬e��п�=6s1\o4�H]�{��V�<�6��;!��;'�����S렃W��-�da@��}�Wᓜ*\=q[Z�
&��>_���F���(Tu���Eus�1��̘Q�=A��Z.����m 4d����m��]]��
Ζ\���,�_{���j�< �&��r������}��,��n&�U{�`I?j�]f�j�x��E<���7��g$����!}L͉{�D�Ap�Cb��.��q��?.�$wS�r�+�[�5�=�?M���Qf4�&���=:6.#�1�,f�s��fU����+�c���0 ?o]�_x�K:�^�̰�uW斌�"�� �o�	1�+N׎��#V�d7ٹ2�bg�տ���vN�%b��x�&��,u"��|�큘.�)��Xi�T�؈�� �[ʲf�,��#���m�~ŉR�YFM�+�O=U��s��Yo�����5I�	��'lL�v=.(�"o��<1*k���	��0K�q�z[��$��CdH��-�>{��.	uE��׸Ft�)�
7�ލ3j��E_��^�\Aԃ�f�~�����ބ�K��'{��3M�5&c�S����Άd��l�󒪐�kZT���-4�&#�YNG��õ�#s���+�x=�u���0�1b�AUE�uP�JyZ>D�y���g2x�$D�Y:����7NhF�ۊ(�šI��+�� �+�p�$(��_8ȸS����)���m����,}u!񸉐��%�.id'���Xqs kDVjG{%�N?�l�)��a��-���yM��gVƁp4	�g�0��.�A)͵���KN�J2��tN��K��7�7Ϣ�/�����hKǝ��q>^q���Q�"�Є��7)�LR"o��q����v!����`�E1�j��Fs���U����[�y���ݵ�S���挡���9�%Q�>�
-�]��:f�d��W����z�q8�`w:�D�2�th�2
�.n�C��d���axa&X��LT��<�� Ӈm,���p�N\���5����X��`��,4f}Ô�j��C�L�B��	{]�W���Z��B+�s�-
��I%��(����p�^�i�}���"��r�]S�૑U�����L��@;X4�AY�%<Ƣ1y���ģe����A��wy;��B�v� c%f���߯��?ê0� �c�L��PPsG�=�>۱�d�Ðy�ʊ*���G�� &hJ��e9��ē�j������"EC�]���=s�D�uЯp�����p|F�!���u4�0�7�����;3$w��!���d3���{�y1]k�"X�P��(�4I�_�J�RD��^+��(�cY��[�Y]L���F�f~�6� 1�3\�%(���cj��@�
>]�N�k�4W�k�sA���"�`x�J*ޅ�u+7��oK$ƋX`m��pmk� L;��7���w9~`���$�XkA!�Q׻�#ۨ%�J�HT���Y8GAC���꿣a6o�o�,����w�j�O���v������"t���}W2�m_�H8�۔�x@�_��R��%Ǩ2�S,s"���J�>9�v�&f�S@�e���o~(G�<�.I��v�W(���с�$E�����“%)5�������v��ݲrx+��㇧��`�ѐ�*�YVJ��E[ǌ�,fo0R5%LY���F6��+��lB�(������myO�{9�L��1��(���ƂyH�5������3M�/�6G_��N�#��=�1��jaYd/H:�k(B=x�$E����Y왲S;���Pz�9��bA$�����K���rI��U,����#�`^0�s�ggJ�XN��l=c"G��xN{��x�ec������:[��v�~�?�pn��>!z��i��� ��޽��3�RI(�$�����c):�������ˤ�{m���h�^� ���.�q�iv�v�3b~���сIvK�m��h�D9�H�G�_!�n:9{����7I݃!�8'��kb>6�LF�y��g�j��쟤\z�%������6NH�{7�Ɉʀ��	)��c=��^����<T�׷8�=}�k0���m�|?�w��_�۲D0ǝ��p�Y���e#0Is���f�g����yr�_[�����\��)��&wA��	Mupv�������;T�Q�(
/&�戫�t�����D���ȉB;�	���i��9��/��%PR��1yo>.�;)��ç�ij��X.�HQ���Vf;�!�0H
�c�.3"}J�[��*�<�vʃ7a�^)"d��k�����⫷���K*�ZaDC�BV�E�������x��3e�J�:�MwƀRW�6���܁�Z�QĢ$z��>v��ݢ�d�b@����fb��&���[���I���m�t/7�+��m��e��O��I"쐕x�w���=4��[u��L���Ce�b�����lwՖ�N���S��z!�v�9s�-�UT�?�y�0�ni�I�E�|�>o�[�Uh��Ǚ3�q���m4�6����
4Z�\����Rk��h�EN�����1t2�Eˇ!o��9<J��q�T�Q��f2�D����/��1�f�J�����;���;����+/��EJ�����m�P�ۆ�����~Aė����_�P�Ca�]�/T�|$}z����,�-H&g�:5�Xt��d���ܘ�qe_��{�l�!O&8�[*��-!��	��N�D�ݘ�b`��/��e���N{���Fw�uf�P��!V�P E/s���Y>�+`��|Lؐ�t���#DI�M4 _��K76��@�2�6D�'x�ȳ)W�h�A���Xm?�\l�_��Cs�"e���8	Q�!��q��J��[�V$�4�RX�*Om`�X���4ysL(���w��Y^YΦ�* ���ݭ��,����x�6�7�&����1FJɎ���˩�c�U�lNc6�_��Q7�b�ő|H�vexi�<h���;����T#ѕ�����Gwk.P����*��C�ws}l�?�l���zkA�0$�d�����2�@L� aM:�3�z�g�,��m�x��.����Czt�y|H= ��˷ʉ�������d�=���e��i�;�;��g��n�E�W�<3tEh�I����N26�5b�����Fڬ�����/r�w@�����r�eoH�����v�NSw��UAR`��^�����A\���=X��
��e�)��)ڀ�'N��7�4�E���/���T{ʉb�;d��]x��϶g[��JΈ���O�5���[_��E�V�*wY��eJ����3���K��&Wg������f}�byJ��WB��r*���ۈߋ�bB�B��λR: �Ȣ������9�%s���������i��ȩ�O�$-��a���wY,�ta1�սSC�㾦�S؂v�3\OΗ�L=qD�V�P
�`>����n��'�J�c1��� /�3F�	.h�'Cy��"���A`�A���OR����V^?S#����+�a̓���N� ����������F�@pV�����D�t�1�AtF������_��A������~�`/uÜULa*G�X~�v��"84hJ�6uZ����{Z�Nİt/�����h�9$��N���:�\�Ƹ�A$�59p�~���hm"���9FSm�h��;���]ƾ�j��Jv2�e���<>R�2�[	}-X�����v����Fle��E�+X����[5a�eb���UZ�R�O�84�M�	�r��x�����2�P�}}G�+�yxu#e?�>3_4����W_�$�V�y������oi^�q��XV�{R�h��Cx��PӹZ(��X"���fB	z��i]ш<"b��h���kM�r��?�9�_%5[2ϋ%ϦH�w�آ���QD>!��sC*߮=oA�6�[����P���
W�'=��@��~N3#��5euLG�E����5��\��y�㲂!SU$�M��
�����Qh�T�6�����11����Z�P��3~��b����T!�rr��NL�c�.�W��]��ơj�$���l�M���[�R���N�J=�q�VBq���K��~;` �9��W�`d���<�����q��'Aq1O�t�K�)�����"rZT��z�f�|�@�<ل�O����,�?��hx�K
0n	�m[{���W�X�����1!��2�x��q��f�_U�kV���`�607�u�0�b� %Y��T����D�@ܔduֵcf�����Vּ���b�wot��)����~�*��YBh��{�]gg�|�&�=�s�0Y��X��Kr���JC��[�O���򃖉�%R����3��麗J��7ޙ�H4cu�F|u��'�bL��3\���AGŒ@E ��i�g��.���S��/Ki0r�o�[P�����:���R���5av���`�=w{��~�O �y.��ԥ��/N��^���ӡ��v�E��o�u��<R�:��Sr�c��� �5�5��p���L�����ڱ���� 9S(E�K����ZE@�Z�z�_�]����Ej�֑�9�r���~������g�	{�B��i�Ƿ�����A}p֦��ጟ��m{����q�%ѓڤHXJ/���h�<��*	�l.糖H��i��ֺ.��=iZ�T}*�=�2M��e�R ��x�.�o���C�(�A��z	?yP~��2����>-�嚙�}�6�v�� z.=��z�N2���z�����[�xH���A�e�A�	����[�ݿI�r��0ˉ"T��L0�.�h���ش�>&��HpB��U�,g���4�A!2�\\X�ŘW1q.h}F��!)I*|@^pو����ٓ�n��݁�z�!�-���WH�?���w���2Yx��.�#��f3&Zy��0�&�މ~��
��e �Y@ׄS�0����G�|�o�f��$�2kY*�9/�@KO��7���zC��I�-L�X�+s{��ev ��_��6fɏ�u�����?��O�de8N����.����Լ�b�s����{*��*]���l����p�X�;%⹄v��W�!�
��$Est�V����$�4l�RYN�9����*�R�� ���<[�!o罼���+tƿ�����ѣF���GaƄ-a}Q��@�OF$Uh����������ɤ�q�����c�~�{��X�Dc��}��FFv��x�h�4\��U-��I�bSrAf�v�_f�U�Sx $wY9�������E�W��� Z"'?']�]���W�mՑ��W7���'�se�wR/6��]-��d�ZF]��'~_�i#��Nʌ<�y�Wnr�rT�����$��s�c���dWcD��l�ca!ݜ�T=����#��]�S�_�!�7t蓞�����˅|������_�v���� ��7��芋�zB@����v�t_:ki��bO�Ӵ�]\�/�aP��xN&B?�bB���mQvq��{�@�_�4@��.��a��
T<���>|_y��'|���p�������3����?Ne�/3\��J
� :��%aY�,WK�)|M�����[Ǌb �{[W*/K��2�P[���s�k��Ř���k]x��KI����ۛt�X�`+�xȽ�z /�Q9kk�/���Q�/��"��>��uA�=�g���$������b�s��0��P`�*1�5����(>d�.�$��ig�w����`�)����b�gm�d���";��17��e� ?
oUl��r�,۷�q�	c̀ԩ+g���>Reb���������m��S8	�3+��q :��,��b#��z3�~j_�Q\�~��x�'�L����Fyy�87w�'�7�`�p��x������Xt�{R���ۻ�����n��@a���D@�k̗�D�ӘQ)�_HT �S!|�50��dȾS�#܊A�%�W��w�x|�R�.�)��^Gg�Z�f��;j�iϹaP_�Q� ���P�����#|#��Y����|V��tK}%׀���9�m�Ӗ�����_K��jc��R���?ơ�:\�}�%[���ƩV���7 �k��k�#If���Ҩ8���������I����D�;.���`�2��z�r�M��9����S%
�rӼ0�&���N%�ȶ����7��/���,�l=�	zNREͷ@�,2�����׏��t�
���DC�>	�nuFrH��bVh4�]��g��������, �B�.~�7���/��� �{�߳�X��c���fs�i�9+��\/����ލT(�O�;F!Ϙ{�m�! ��8ih����D��@̄�5}Y��@�n激���>�H��%׿�n��A��/TY����9�	���l��1���LL����֑d?�Ʈ�X�I*<�Ed@��������.
�;��`9I͛��4	TU҆0���8x7��^_I��4S}��o�m�dm�Q~D堝������T=���w~9���Qf]�ӯ�1gW���»�3��6�i5�:��pZΓ�ut(���G ��y�8Dz���v��B%=�P�{z�(]ħ_���bݳ�c�����O�ϱ�x#
�97�6�P���.�a=���K֔e_\�5�;  ����/�l�3��^|
��6��!��2�����>}g�q�r�����쳢��[����fCeD\l�"�����N>��D�c����*Fɪ�!4#���(w��d�J�u�zQ�C:ej1 ��ke��&���_�G��_ ��빗@%Z���š���2ؾ�2A�?bP�=�9E��kZ�U���ěn��N�� �t{��֩��B%8q�O��F��X:*�W6B>[��fٟ�����߾U�뾹��f>���N>����hD������s�|�B��:Ue�tθ�i���c����PSV�X�C$g��=�O;x�-�B�_�؏hl� �צj��;9��Ȩ��d-��h@y��z��\3XoHy׺Qv�J�����SК=�mhS��^ ����DA�C�\��)�)���e�����E�!*� x���#�=17���{:�a����.��{�>��F�	w��&b��r���0��0�lY� ޻uH���Œ➝㾋��-���	}�󂡛iK"�����������|.�2mP����k`)�)U"Op���ST+���Cz��L](#���Z��3�ᇅX��S�G?�t5*������j�J��}^?�bl�et���҆��	H�ũ���M�i��U��4�݋�ǚ�n��v��"4�5*t;�I"�f�$HF
ު��U��2G�`���EVyO�+\ť�|�2U]�h�?�	OR��_�����n9;�&=/�9ށ(gi{����o�D	�&�j��Qr�����Z�����^(����b/��$��<z(�9�T��>>0�{.z���p�����vjߚW�+�P5hQ�n�L9�?��̃��=7���W�ՁX�/̭b��kv�0r	&�1k�LZ4ڛ�u���_=�E\u[�+Q��OOG��|y%Y�x^��2;�^yM���O$��}����*��:�d�#���!���\�p�{�jA-2RT�iػ���,&��-�7}��Lc�j�ys�P�I���
��T�('���x�Ӳ�^
^R�)e����;��.h�~�����p��Y<�yŁeн��(�P�qҘ�+nS}��ꠎ�I =JzG8��%~^�.+�0߁�8G�]б������ׅ��ʈ�2�sr�/R ���B��q�ω�7*�E����̬�@��/�zy���Ò�p����R�Q��W5�`m��QZA&J���;�yg�~�$?�N>"��m@���N;�5pq���^=�%v��.��N��^������Y�
�#!eR��_���0�7tZK����W�bf�~���sKj��=q�1\C��I�B�Ì:�N��<L"��]���/�#ǁbA���1F�v0��,ݪ�)�m�fr�������o�9CS 2��Y��$H���83%�2TϮ�8lz�p.��0 E@�E�H�y� �sT[�����M[o��1��ʈ�M*	_Q�����R�i�|0�ܛ�;���	ގ��s/`Bc���,���z"�C��uV���>~�Y�zN��O����^��"h��o�.-���TP�}�F�W0��D6�S>��o1�%�L�5��'*���B�Y��k�ȱA*���]��=��2@7����+q�������A/���f���&�}�v!��� xH�jHfFÜ$�G���h�S�{�v�m��x#�Q-�f{8�Tȫ�	�{�MM|�{����b	�]�1�..�md��E�{�`�ð�[���UN������j�J�J�j��*
��~-*	��K�����zp�r]����M孲�KryAp?Z��Bv!sэ]��1�#�ʍ�&!�/e;u#M��RZݹ�@*�c��덽�[,cj0FL�|�<rt��b;bJ���;�{/�[�=��3O�CAL�5��XvO�U��l�<��Ht��/wQ�!`)�� � ��^󹎶����)����:�z4t?]�A(�_��!�|]����[�
K����(L���ao�)�{�xcǪ;d�ǆpQ��Yè`��R�cuf�(%���1%�=�Չ/�����p>�m6/����*,���$07iD��f��VO�k��>�����ҧޗg�B�i�<
��j{�"��)U�p@���6�1���o�6��t��`� *S�0]RO�g�.L�|�A�#ـUq�M��
]�5qhwɌ��ʆ�l�t���m,>�������2����is���"fkâ��r���E�)�#1Z4��L���OW3m �NC��s�e�a�7+���Z��x�+Q�(��M.a�D����T�L^��կܳ����;*_��sg6er�DT�`����~nTJ^�EI��5jVE��_�R/}ă-�j!��{1���'�C����@{hq\+v >�-����#��ZG� ��y�{��"و����qo�QF��y����vw�|)=r��hH�r���>=0}�Ȇ4����Q�w/�Hڰ��+T>�<Ng��+K�8Ow���1^Z�f��������ԑO}�CN�AR̀,�]?;�7�2�m�L+jY�	?êu���~�Mj'5~X�S	����M�:��֒
GE����#�:ґe�D���K5�i�Q���3���� mvI����_Ê� ���"�o$y���PD���A�2�	>AcC���֏֎B���e�>@&��ҩ\6�>�*��es�5f0C�������������w&F�^�F,\_$�!�?KZC���O�|�a�(o��f��5�����V��W�������dkj�0�n7Ԥ5���	D���X8�Uk��;��B���vWSw$�!�a��%,��(���������xk�꧴�M���4z��^�v�pK��|��#�;GJ�ʗl4E~+�S���m[$���6<�BsPTUG�0���Y��W؄�q-�B����֯�w<ސ2��^�_R՛I�t�ި��ʌ꧱��-Rz�]����_�FF8��� *��L��Og�\��U���I/�ɳJA/�X�?�,\�ud	]ݚ5H�q���TP���u�
��d�@�h�#�
ߦ;��i� �l�rtR��R�1Ay�F�P*a�ݸ����֋֪��zs�)#�F,%��=�`��-�=�C&�����y�?�"�y�	�n"O^��τ�l�9S�P�6z&7!���#�$'���ϵ��z���^�Xc�u�(	Lj����0c�]�jn��C�9����6���N�xI<�k���W[g����ˏ��PK�|渓������2|�woN�������w�"곫{D��!ߐ�fGZ!�G[!�1Y��Ȉ!톻�|�'�c��[.�9�`~ǌ�N,�b��Z��R��(v�$u�HXthw�Q���|�x3X�bk�.璲�2��&}
��8��!(����Ń�V��[��q ��{��{�8ךn�����+1�L���]f���1r��{���8|�p$�����ب�y���A�M6���
%M�/g�qr��>�zU.�՛�^׹�򎿱��ug�i��I9T�G<Y"e��bow2Q�����'^���� m�AT"� Ew��0�a��h��y�X�P�vb�
`h͎��5�չq��f��ٲ�3a;���гuq�Uڶ��r����j�� ����9�������2ٰ����%�Yjlof�e.펵�u��i�0�}7'n�d��8�\���N�� �Q�	�L�j@����2jwz�G;�M�OJ�����1625Y�g'�v#�=$�����4��4�q,AT�\C�0�zwe
g���dJ�~���i�O����/B�Cw�S���	c~�3M�u`fD��E3/���Ӿ���U��a���
6շ��1\��yH$����$rAn�!q�8� Y	f5�t(+��6��׾a=/dN?D 1B�x��'X����Ź�0@��@6��r��f-��,ʍ��L:�b�ap�\Қ^	�ءbd�	���F�w�(�狧ڧ��=�������guNZ�K���xx��޿�Gd!��,��:ɏ� r(/Ш1�K28#�Fl ��Mß�L��1roӜ�(�(���I�P���A���������N�"�&�
�` �9�o���*���=�.��K�&z��5��E4� ��]t��35������r;ɬ�D*%�������qxKϊn��D�{U��#����A.V�U�J�I)�<�х�����lTv5�Y{˕"�G��1���X���}�p���W� ||��&����8���).�h�C�����Z+�1[�~�%Ki<Q���<m�iHD �Ѫ��@I!o�ut�v0����nG:
��m�x�����Lp�!���D��n0�'���N`�I��)���O�^ċп��e"��{]]�U��-y0���n�=�<��gW) k/-�Q�����<z�� ��=x�~�_��{���T�>�K�u`N���J�������%�L>j����q�>�M�Ւ��^�9SA�^��qf8�@1���0О@�����vgë�8�2��I�����q0��&�,���j����0����;MY*3�v�M�;��j�c�/��6��j��7b��D���h(���&�d���.�)!����_�3��
�Z��U���'U(�������&��&�n2&<������_s��ը���B_��Q2�v{�|	<Y,{o�P􎑣d^OC,�`���,j�KK���D�2���$/�s�S����
^�����$����[�tI��/�k&Ev�����W�?^���٬(/9>=�e�qS�:'�}ʫ"1�v�{�����+�`υ��]���)zy>��m-��G6��^IX�SC�ĩ�ֺ�#!��e��2�S�+�<�<ʳP{&]OV�K��A,����=evb�X������E����KGbƷ�z���E D��8Y�/]@�MT�
���y/ֻ�^1��s���`�h��Ёef%%���X��+���[�~����x�)��`c%$�5Ni����>t����-����Tߔ0m[��B�c�&uV;EĈj�)تVjCj���|.γ�߾��7�԰9@@�Ѐ�!������q�Q��F5e�]�K�})���c/35�%Dm��=U=r��L7�w	VE���L��p�3|4y��y+=�:����m^-tu=�.E����>�F�4Qr��u�^�����IL4v6R4)� ��Z�m(y�Lu�T��0ф��E�íG�o�}�����UË́]N�kO�g�	|�����&��T�^�g� ����:�O�[�:����C�uw"�V�Cf�L��A����){���F��{�WM��(�.��u��u�{x��wL�s�f(j�����Y��td�c-�ģhP8Ódi����W���m�,ɹ	S^��jQ�u�1G٧��ŭ%=t�ٝ�6�q�,#��eA�B��L!�������(��	��P�����ek��	���;M�V�|w�BS�=l�PX�nr���_"�N�U�b���d�i��5o��p\�ʅ����碷�t��i
 3×j�C���WNP�$�$G��7���<-��Z�_+��ӯ�&J�X�V)i�I#���R
���Sѷ�������&Y��P��)�n#���ְ2���ϒ�R/���2ӕ��Z�6�����1B6R*���$��OR������+�NuP,�F���}����0HݏR�mC9|���,���f#�\����;���0N����xN��Z��ϯ�F�GjmRR�nG]���-9�>C��1������ڧ�A�h�>�ݝWa�y\k Ф#^/.�^P�T9ս�����g@�Y�:mE\���㏫�%�g}�@F�������<�C�o��<r@���v]�!��~'(�����ζ�4.@�^��[�ۥO����J�GO�_\B��K�@	�����se� r�KA;K<ȡ�'w.�rb��pD��5����&������+���H%V��; 5�c[���/�ޡ�V��BܰI��2)��z00��'�‬�1S��W�q�*q�*�)�9ֻEMt���o�hf����'�����΁Hwt���m�ʞ���.�k��N��K�w�%��[g�v�{�N��.��	!{���%�V��9��Wc��&��(6����t�����f�S�{I��>�"����M��ZU�G},�EN���N�*F��>����Ad1:�5��^T�SEu�뗪�������@¦�TS:��Z���f����i��<��mvHʔ��<��=D$��p�w��Ó;���4ؾ�q��8I�g��C�^���[�C8�2��7m�c���Y�U�z ��y��RhhX}B�^U���Z4���yT��׀����J}9tv��{y��>L���)r��[�g���tT�
���"K��R��O��끂M,�X,�H�r��/��(��P+��U�$��mo0U~o!�B�&7 T�Ҟ��ۼyR�}@�Q��d�~6�����e�h���$�_-^i���lu9�������f�N�ŷڤ����wk~2`���ܴNHU��R��`��w�թ���ų��ïٻ�޸YЋ�#�#߫��n��O�8���.�IW�&���n���*�$gщ���Wg�5Q3H�:�ٞ!�忦�l�<��ܢUK��i)?��,��O���_����B��n��H��D"�̶\R3�6gƛ��؞!E-��Os�0�HL��;x9!����Q�>�`Uݛ�GR�(<w���������3%28�^J���c�����DB����,���W:#>i��8-c$RT�.�%ʟ�9�����@��^[.˔�	%d�O�f<�T�W/��#^U��H��$x7[�J�7!޾�rQ�a�x������\��*����ql!1q�QK)-�Н�MX�\o�*��#lQ��_�'kH�Oܟr�/}[z�l���12�^|�x�����tw�E!���4��i�����=p�w0Z��e���}Z�?8f9F�1h����Fi��~����*��8)#�rD̉���>�jI�UЍhy9J%N�\� �����L.|�lĺ|w{�+�o���� �9��d��P;�~F�4�E7�l����?^�tw�6���8��+����z�#O��C>V�W+J](��"=����/ �㺊<OI� �Ro�+��/?gA�ŧ��s��0y��謎��HS�ᩛ.��h`Q�/	%��N�������K�*#�ٓuV�,���@�`�uo��;��W�2��!�1�l�j*Gz�5���_Ũ��"�<Âf|Ӵ�C�W�^����&��L|��i&R���݃��,��-����Zi���IK+�:��%9�%�?iH����o��;�K��q`*����&jts�y��v�L���.��<�m�8Pᠵ�N��߮Ū�_��M���a�?�IeA�5��\Y��!Rrg�`�#K��`cf��9˃�dO%U{`b�>�|7O�)Ͽ�ݙ:bh����#�m�%����k~@4S��j����;�G!@���	���.i���t�~t�?�qL�tz�#CE�� �H:oV�8�fC����ʞ�L���������v:cf\��7���p.R���a�ƫ�}~��1"�^{{��`I��׹�#߫�sC���(���!�����'��h$& *Pz�U"(;���G�
�(o�Q� ts�9�'^pN���נgh�j��)X��c���j�7��0c���v��-9TP�+,���4k`�C�/�Q�V�D��j&!9[��0���Cۨ���7*�c�A��p+L�����]D��c8�<6���9��<��r0,��s�ixU>� 湌��iu��cBq�ؔs{ō��u�Ch~�Z_�I��p��v�Ct�(Bz�nZ�b7m��k�aƹ�:����5�h�G����A�?N�N"p,̻�����؟�n���+����7�o�MK5`�0�:�oxn�uϗ�E��u�E���
?���a9�{�>�s��X�Lp�`3By�+��)�ps���Rp�QI~1w�؀���F��f"��@�}Zg*�]�i yqHy��: ����Ѻ:Ǿ��^��xt�dP���m�EsГeX�@M,)����k4Y��XIz�L8�yl
O����];2o�b��}�ܦQ��24x����:�7�P	 8ӂ�=z�,Mtjx{����	#�&��`�3R:	m��Q�艽�⮱=�_o����~��X��]�a V����^��ƴ�k���Ő1��-}!�mw�%�C��b��'�ׁY��X@X'��=}L\��=���Ǳ�l�u�ο=�E���p��6[�����槜��@����Alyk�[��j��Ֆ���dF2QV�VEe�Dw�E�O�2�c�/�Cm;�k�֓K-/��	��m_o��Ϋ����U��5)~�ѯo��Ѥ��-lOμQ��1��+�ȏXl_7ʝ[$9UOZ@�y�U��s�?��v�������Ȅ��
�V+���{cUW��̴~�4��҃��_���U��J?���,	�H���J�d�s�s�0
��E��/�� q�B5�����H��\΅��;����s��F�%�:��,ۃ��bk�Kױ�q�O��(�C���yr�B0N�iA��"��̤��p�/�;�ZcB�O3gϨ�9�G�A� h��m��Зg��Xk�rϧ�~��V
@��s��v�h|�˥_��|�=ׁ�pE���ͼ}R"��0��7��6;*��P�b�i��/V��4Ҹ��k�ӻ�q:�ZƠq̗'���Xpv# ��e���w�Ê�����2��<"��'@]�9�AN� �m�Y�M}/D�d����#��j"L�̫����L��*]e������M-}-_fct�<qh��@c5���7~kܾ,�T������9�z+W
ֽ�0�)��Fd�+Y�
B��B��s�;�N!<eo�.S���..,���\%�^���w����ɫ�H�ڠ<[R�n�����}�/�U̷�.U0�o������a��oK�dml�@"*,�cL�P}�1��
?Jo|J�R�«d�N禀���D��$��q~�����LRk�����f����)-����lf��(9@c#���%1F�$7����Ր9��x!��Dfn]������˘KsQ��))�+ׇ�f�[.c�~�n�_!�1�y���CG�ے�G�{w�OI/@��t�f;g�}m�jP��	+�&EUh��`��]b9u}m���=Ri����w�i*<�L�E`�%��H��:�t���%f [�(|���U���"[���͎�����T��:�T�SX�RN��6�3��� X�|���?����,��u����O�"ʂjEW����S��Z�vIUQa/�L}\u�a^y	>Oҕ��{�pT�e��V1�ڴri�p�@4�@�O�rw#O�86%܎����>���i$�5+7P G��?u5_3�m+;.mCk�4�)M��f0'J8���R	��j)r/�Oa���hH{���E�(]�?�Q�ie�"_���4����?�Z�":��Ѣө�c�H|�g�s+[���1��c�G<��������b3��Wv��E��H�U"�*���H��܃�4����[~̡��F��=B��yBjb�}��F��*�O5/���� (�
�3�F#9v�~��?,��K!�+&� �12#4\��]ScY��~ڈ�L-���Gixwi�����y1�b�X�}L��i4����
m�r�e?��+���|H�r7w�32�̉�p?xa.�q�w�i��׬!{[>�o�2w.�,ϒ����m��dj����+_j��dLyC<����P�����C՜��K\����ކ��'����CN��BZ6G���3�&�Z��O3y���3p�TW����I�b*-NJ��x�R��a�za�n��f���n��9:c�.�mޒ�|yb^B��=����Bc�zw2�,������I�h�lg�H�����̭dM�dM�(hϋ~�Ԣ.����k�����|dd[��oE=�I�F@���+�c`偝�m�c�� ��TRЛT��H0&諎���{s"l�])ɀ������Tb�^#��beKi�f՞��FZ�F�"KK�)�LJ�U)���wx�|��2ez�+.}@�:h� DiD�.�7Q�f��</���*$s���3��6}; ��~%�i���s�"l�,��5ټ��q,6��|H�������r~8�..�ja�J��?H�"8��0!��ts���n���Sz��J����B�NJ>V�,w��L�S  =�c`  �������5��(L�$�/����	,��@D��	l���댾���}�H��$��Q �^��|�;GزA�]H���f≙����}�3�_�Un�,pe��Ԧ����GK0�A��Z���X
�������퍔6�2�F��~�Ң���>��Pf�|�AY���L�yj5��N �X�O�~O$�* &Ǜ����q|����� ��縦"�P�?��0��5����4�T7�u�"^EIJu���RS��3��w0*6���V{x�+��pe>Ja�\�"4��k^����`.X��#�h�ɚ��㒍�nk"U��I���)-��v��5���è�f���?��f�q�����XR�YɌ	�����>����
�C9$j�@����O)�������NPڑ9����c_)�n���V�(ȰI��	��JB���A������5V�T|�h��,�h�U��G�(�p�`̡(�u��X믓����탍B��얃=����@U+���������!~������^g�a�Y-�3��K�K,��GNy�^}���Zǀk�����X��F=BW��L����?��O�J�G��s�V��,�LS�����i:M�����ʴe�F�~�o�q��$ë�����|��9�|ڝ�WlK� �����e���-�,r 	��� &�!�Vx���M׆��ve�!3�`�9�O�4�(�#��T����Z���-X�;lH��v�6J�0d ��@�0Fbm�f��t�w�z��u'�rAI~�� Gd�r`���>�<�\];��d��)T�4�'rp^0���]�U�Wk�(�F�%4]h�\j0����`1�L,�	�-�}����xR���a`q�#�G�*2A���4�V�`CD`q��@94)�X�����O���1J0�/���ꗒ��7�D����J�(�'Y;rH����b�r�؏2��&�x�fz_�/2�[�ʄ��.&���d�q�m�{F�ѮQ�'w�\9	-�೚��y=Tՙv��oU<(�89���d���zb6Y�����ǒ2�n���&��	~ʲ!x��C�C��jO��-�tL��Z���\�a�@ĴJ���S���B\X`�E$�5������Ҽ�M�(���W[W���U`��MՀ햁�G�?xU5qH����栆4X��Iv�^D�9;���V�K�(�tm�lm�	��M���p�2�$X��^�D�%���D�;�3�s�f7�&'A�@���>� ^Z!E\��Z��p_v�鲳w�c�9̚-�OL}^O!�������ГӄN���fǞ�@-��.�����֝#�ԄZ"%O,ǵf�*?�/����t��0��nV�XL�}�>"� ���Vhk���v��x)11/��q����4�,�D]�~Gd �&�pzHZ<�gEC#�:�)Sz��c�3�m�;C}
���A��(�B��9��^��Qj�yU�J̨�x�D�o�N�NU1#�)��ES��d�A}QR�t�k3�G��c�������E�g8��s�������A}�!Ş�+Zs�^�`�V
}IWMs�b:]d�+~2N�RX����%<���5^Z�x_�����v��,�/b�c�v���/�o�6�]�X���/�D��H.�R��ۧ^R@�L��
��4�p���Oᚙ9�GuyK�4��l\&ʭ�Z'wRVu4��ׁx�[�{��4�k2fM��}�}-���M���������5����L z4?U%�@򚂫��m�z�5�K"J���J���qH��/�='k�9�D��[h����|D̩T������/r7���p��;u�bjǎ�j�ü`�\���� �_�j�åC��n�~�q��	�5�u#��D)�j_�h�\��cu���X�+]X^�Ok=+�B�(��r�*�]�"��S݂#���v������w�c���bX�#vf pH����+u��_���ѥ7�ւ�A��i��ۯP�7�*��
��`�&��	�30���XG�������WX�����_-"�������$@�o��!�S*!��&(�����MF�X j���d�甽��*D�Lc�\���	BD ��r�N1����8�^����v��'�g����3!� P���(�pU��b��X����ke;1�< Y�����^�c���sέ�/�(3��Z���z�f2_g��!�O}"�+��T���k+s5�g�	��W3Y��;}��i�|Q/�/���XL~Z��3A[�[Bh���Qu�7��DQ
�؟��,�~�E�@�vz�ؠe�L�ۭ�ݫ�Rؿ���uE$L�\�W\�[���4=a|���x���3�VC��L� ��KD�d>6�"��}�j��9џɘ�������f}�Z�_1���:%��������Qr���RyK�%n+�8[mUz /l���g�Oc����FS���t�-��y�D�qc�1HjǾ ��dH�e�cֲ��E��F��[�M��ͅ�-a����ÒP���`����gA&a���C�Ϲ^���|l�\6��?S��P()��� ��Q.��IY�<��g;��s�Ǡ%��
-���W�6�kn���?4,�O~�\G�)nl��JҞ� z���	�Y��Ӻ��	C����Q�&r?EFl�:rƗ�}��;=5��E�~�y��8L������$��< ��	��O/O��P���Y��Jz�~��a�	��A��U�ϟw��X���K���ZD;u^V�m���a������Dr*�vr�F�[���L]�PX�xr�߸�d>U­��2 �a���w���W7+��MDu����z����6��Ʋq}`'�.��ƀцa2t4j{���Cz�i� �BE�/i��7�M�u�:Z|_��s��4K��9^�.� ���G�|b9�����u�Y	V}���Xl���v��q΍���3��� +�d�� 7��F�@9�N=��
����3�ܼ���p�ˬI\ؔ�YԺt�� X6󃭶^�ب���?���Cx���)�BZadPy�z�+x�̃�U���|�O�W���KJ�տ����PhDn/C32�=ME���&�+�AC���F0�T��^�:
1����V��*;�?�\�ҏ�s,yk3�n)v�j/���3����_�&��Δ��.P����I�^��`�U������A&E��q�i�cv⸜&��_��T!�,��*
3N}�|,�1��@g7�<߂��d��8��ȋI�ؑNЊ�
�(GWWq3�h�"�h�/	�|/x�Q'��ma"G,�fY�1`9�e����Q(�O/��7ڭ�T~#@ߩٻk<��g��4Mĺ�)ڨ�a�=�{���R�\[l�6^��7��
 ,���<6^�΄�$�1,�0�Gfxc8��̂nC<+vJ�K�OzM���=!aۘ!S%�q�pb.$I6y��m�v~����/;[�+�E���oF�iR"��8_��.��q��zL+��r3����C�ȋ�h�.���"41� ?�v�0�{��YӐ���A߰���H���o�;� Ӟ��n����v��?���&���x�m�P�X!^e`{�R�V�(5T��(�>,!TМ0	��d��GK���6̭w��Z�y�lp�"�;��A{H�a�O�&ނ��Ƒv�P���6�\{�Wxbӫ�u�H�*V�p"hJM&f�ѭ���/�J�HQ*�"W�����ʭ暘���(�VƳ:6yڳ���g��8�4�$b�I�g,G��zC
���� E��f_����Jd��B�a�qF����[�y�{�^$�:u���i5�Qʩ�%���+�q�W��<Kw�/>��<��:�����"�3G��c"��q8|ASvӏ ��/�����VhH����[�< �7�nR�_wC5K`<�U�=4��j�.�kc�'j�~¼���u���:���ȸ�e>�5�[DB�68���� ��	���Rg�g��>A�Ο��x��x(�Oߋx�F��ط��u] ���mvH^[�O�'����3��R�yf�ΔM�Jv�7����IyB��b��$cE��% s������H:�f�0�����gQ�b�a8�zt��.sB�������#��K}(�����_�I��i�s:D���2�"o��Q!:��Z�m�5���n0�K��� t�<�A���a=�=�#�-�,�]���@s�K��K®Su�x?�<��5q�Q�zP�(G�'�F��X�|������ƺ�M�@�/푗y׆��ϖOg��t��B ��F^D��^��:uɶOI����b�5{�u�_,:;�D�i�k�E'A�)�yC�օ����g�����-� �B�9,E�������O
e@�V@�h�_Za�r�Ë�*[<��"	x���/���-��w�k��\��r�6�6�ftf�(��v���Dj��+���[�u�:�<W��7a���L$��Sh�ȿ���l 	�ܽ+��H���Bb$���]��1dLB�G:;�Wir��@ͻ� ��|r��P�P�5��R�軣�ŨU�5��g*w�uO��k�{٩x>��(m>9 eS��a���U��P�LWE�N���Y11���d�mEVv�7@E�t��bη��&/v-axw��OR�F9��w7�6hʹ�:��'v;�C�ְ����
��E�A��9d��u-����;�(/7���R1��¹Q1|���ܜ��/����t��aĩ� �E��Zy�N�z�L���/�A
�/���J�_�n �a|�<�֋�Q"-m�o<��j���<�zv�v���@	!��i'Է�k�*q����7��8��o�1zV�9`�V�E
G�&�-��]Ǧ����aR5�Zr
b�F�nF�;������2��
�9)H^�H���D�[g��Qa��=eI�~q��eQ�Ǐ�XP/���d�݌���!��2�`�!U!���P�y�j��d�ȢH�5�ܤ4���z��x�
s���=$^�L$�s�+�[kd��sѬ)}a� C#0�z,��PF5�p���u���B�d`��G���,���Pe��mKϼ��L&ع�u��j�q�di�#0 ����W�հ��}"3>X�c��3�K#�����&?=�T��@�vx��Hy�ɈⱸF��*<@��jvQ���<��ovL���>��9��i�M�hۡ
G&O����F%�	vY�� ���g����q���Ӣ(�7D�e�ͳ��קI>�Eʴ�|cJ�������4�</֕�����z"�E�j[��9��	��5�mdp�¬͘Q�7XT�MH�m2�`�ޟ�\I!��ƃ/�sMG{:u����wS3v��q_���\Y9�gG�28�hX�D^����Ӣ r��F�rl�/�j=�7	�-5�e@���̸��*���[Y?�A���_%b�;�{Vܙ�闢U�N��s��U������󁏎���k�d���2�q�?�� �=�+��[��I=ޙ/'|�� �7R#c��=C�\f��iB"��̖L�R�[���U������ӶL�E,�U<�Yd)�2��wZW���3�~o�N��C8&y0��K�X� zN���SO�%����+����r�UM �Ko  �^/:�/��e}��i1��A+���Y[*Jߐ�x:=�O�nJ��>m�Yj�������pk~�+é��y�8�?��n{:��$}C��E-AL�{�V�8�a>l퉣.��0�;��:SC�؊[��,%�4��؇ 	�g��a{" ��S,�&Ō������j+W��vcLf�>0�P�����ə��Sn��Y`�f6ղF���a��o������'o���/�vl�MZ�If[��Ij��'��6�_Q�{w�����"����:s�#1�[��E��R��f�z�WO֝ɤ��f�-��((�bƌ�ؙ�4.�X�����F��̤��?e->rne~���H3�B����eI�'[Z�#+r����M� z�Ca�DG�U��9R�]��>��`�CF
 N��k�69߉���(��%�t^�<��J+��X41=�������r5:���"nK`��B�@��6�΢����2Ea����+�n�&�,��2��u���d[7Y4c�!s�j�W2���C,�c�&5%�~�������Wq��J}Fe7�7H��43��#�K���O׿�BP��"#ߚ�ߜ�J�ڝ��>�%��Z�n�N�A�:��Ѷ�A4o#g��ܕ;�Z�b'�h��}'Ǥ�o��"��7�<V�8֑۔9%Ab.(�6u�!MM@*
��Zۉ.R����ܶ�W�t�|#�� N�����]jE+�*����?�����VI�.WS�Z�~���C�ƒ�\��֦��;D�:&9|���Z�����wg6�������#6���j�8�����PO���H�p�Fs�zb�%��gk0���0Q�O��i U���ݶx��,�q6y��|m�0f� �0B�\>o�]��[Ix�`�qBGJ��53�VLH�T�2���u� �r�e�2�r�����d6�,�V ��P������'��etc��7������@�ht� ��'�Ւ�`��9�Ϝ�_R��s���R)�ڪP�Q���ya1��C�$o��%2����=-����_�w�� pQ���PB0Ə���`��>�Q��a� ����58����Y~�����~7�D�x���f�
��G+��G�[�!K�a&��`5qѬ>C�G����M����b��I���D�~�K!��4�iQ���6lυ��$�֋K��^n2���k�,%��� \ƅ��}�BC�mӸ*w��sP(rQ��Ӷy�J�cz���0T�Ƙ���tx����>�������(u"�����hu� =�{$�ek��q(@yQ�����$�PŪ� ��������hJ�ć1\�@s��ʸ���'�SH�od�f��Bsr�i�(	jun_:H[W������e����A�i�{����6,���=w>K�֕�r%�C��&#>�K��4>�[��������XQ��iī�<52��]��3��Nqk��υ��9�e��Z$l�O���z�i��S����.W�ב0BE��5��z���;�;ͨ��H��6�(r
���N6�:��_���4�+c���M�\�ą�z6���� ]��	�ᆲ8��@�t�%�I@'�y������+���e:[0�x�ǡ������A"�@�����~Bב����(��N=v�[M��O�|���_K��9��ޝ�h�Ƙ�3Q"����^Oz� }n�I���A&f��Ȕ�i<Pe�����8��E��8�@�P3/�?��:�V'��IV͖QBS��hѵ�Dv��~��bl��x��`�����JDA����~b���f�$���FQ>�;<�9n��$���@���r�MT�J�l�?�ɉO��ө�X�K��デ� �ؿF(L���(�%�b���|�?8�5
��8���1U{ff�Ȓ�|���f���nq`I��ӓ�3'�s�n�:�l��o�>_�b(F�2��x��9��ae��x�<���܆+i]��]%�PG`6��Y!���A*+�y�w��#Sծ�]������x�W^]�Q��I�%�xV�v�#q�^����->�n#�f6r�ͧ甒4U���|?��dH���&�D�Z����
���Om���a�tĺ�Uhk���yȿq�c(�{�^"��C>�K�;� G�\y��*���ݡ�?��Wc^�L�!��vP�����X���O�E�ٜZ���vӴ|}�!3^8���?�Ge-�Gv%�^�\�Z���ى�<֮�D4��%}�v����u<�W2��}��;��=׹����"�lm��Z��yg��#�#ÇjbD�J|J[�=R���M��\K�2�����wA0��H
��C�zE���>�,u����Y�8��)��>'�B%��@PF�Y�<(��|�_�q�O]�_}|���KSA�,�ϯ,��u�B���DL�����#��2q���8��'��t��B�4{7��
#z����Ԁ���t�&w�N,��?ؒ�x�-��z�u�n�� ��[�B �7�G�b���HǦ�wџ*���Y���yNw,Gǡ��J�ID���=�n�0�o�H{����I?�D;*R"��k���ʵ]?i��7'o�Yk-�3�~�O[�������!�b�Ϗ��,4[zu��ց)�"�
��}]u���U�s�*y��o_E�b�k��
j����r��'{��^] ��_�H/��ŦGj>�
h��(�K�w GU���-��8�1V <�j+���� GMV�{����KI5>�6
����.
 �|:s���P�����Bs�{_�G$A�
{�F�RX��l�x���k���d �E�S��A�H�e�W�ȇ�FH+ΖɌKg$I�15���pO#�fISj������t��m�B����GE�/i3���}9�7������e�tl>[��u�͋,��ɬ�LY�m��Z����FP��L��+�q����K�7	T$�� .?�����[��|�eQ�ʉ��j�D������:�b����IjB�YY�2ܓ31�t��*�E$8M����x��
�O*�P��m���N��?P�8֬��K��4���t��>�um�[Ą�K�L�1��۽GY��-E)f�#h��g�����-qm���j.9#��H�W��B��:d��/c�
�P5oE~)���Y{�㩙|qj��_c�Z.4��ź�1��P��쩪n�tK����P��(_7��i�D���:����p�����\	e�-�G���5O�C�
ZQ���[�[t㩤������n
r�Fp��.8
Q�|0���I�!k �����iD5'�Fg����+\{;�O�=�HI]�'"V�|�S�&;�u)0I�F|��k�v�<�g�2H�wq��� 0Y�f|N���L�T{�%��.���bΎv㴡�6	��A5��z��Q�¼��	���P��R�5�ytv�3�V�iF�ך��W�Y`H�6ʄ μ}F�
e+PQ��^�ifG-o]E-+��w>Zkҕ��#��s�X��;$#7�=ų�ǿW�ZF��ޗ��#-
H�P ���j���P\\�m�蒨`<��u�(�u�g���Y��'[ߑ鈻��09�1y�s��;Dʿ�ZɌ��dosXk�A�^V�䙳��4�F����T�V��(N������@��;*�O'fe�������s+�y��Usk��տ��� ����6K4�0o��/ �ʠ	�@�<�KN��\*j�_.����5ln_T�B�(sI���L��A�}�\��'E4<r�N��#'C#D~و�c��ݣ����+��Ta6=En�ټe`@�%�:��e/ŕ��/�����+�3V��O3������?#�-��`,+�ǐHD+���fVi"����8xF7����\)��v�|���o�e��ԃQel���F�1�����;�K�!�z4O�Mz_�3=��$c�F��@�RNB"ѹq�Xa aG����*�z)�4�����t�j�c��.���O�_��C�A̸1$�P|�2 ~f�y,+�>��n����[�@�%^�6{�?*;-�fǱ�YX��k�nR���K�_������sj�g�soM�"�W(�#ysrz��bn?�Q���'��'�z+� ��4Խ� �8oP�um�j��z �R�(������Gx�{jӀ��VG�ӿ%C���H�o���eH?��0Ϯ{�
�`V�Y�JOFZ���ʼTCp��;sȯ�R�_�x�φ�7�;��D��k-�uYh uS�j��%�M?�7K����Jj���F�Μ�q�%���?���� ��R�R�l��춛��Sأ��ܟNZO� ���Ɩq�݃�GQ,H��~�,( z�� �T�([�͔?ݾA2Փvc��<��m�@�/7@AmP-M�_[y����}2C�W�ȑg�b���q��K�>�w��̓d���	�-���G���f�3�~)Q
�[h�I'95�"x�.����Xs�#M-�de(��Zxa	x%~����rf%�B_�����8���Z��Q���0�%ˢ*9�N��U)	���<?�,Ͳ�06җE>��O�Z�< ��sb�� �g|Q���}�kZ*�خD�>�r���?�/��T��[L��n��P�[w��:�.�=�Ԍ�޿B�%12�e�e��A�5Ԑ� �[	�"r%ş{�ym$~Q*�Z�۶#�{k�\�rZ�Y��:1�:
�ɑ�.5��F�ē^�}�W�a��d0�˯6 �J�A.0"� ��t�J��j�!1�BM? 3��K��V�n�o.sJ!����8������f��1������֥�Kx�E-�a�¥�(#��C�(�Z�ӝ|���:cg�哞 ���3 �l`«�f0�Sf5%]�,�M�R+�z����V�y�k�b��& � �؆���/&0�|&�%6�i�u�R�s���r��G�#�� +�#��̜�Gx���B� �[2Rwf��]e��/i �@�	����tC䯖�p�Ȥ0`���!3r�:��FF�_]��D�H@[f�y���$�`�4�v�O��
}s'�ǰ�9Z�9,�i>��$�q����b��)�'�7ɛ<+4�1?@)�pT#o�	���'p�٠#� �ʤ���0
nx�/Y[m���f�S���(�l���r�I� �r(�G='����Q�3�4� Ct;�A&�)/�-&X=�l�t����D~��m:��RD]� �4	��/𷆰ܟU���e.
��~lB\6�534�H�|T��n�E� EX���h�_1�㓖q�oO��Z�K����Z����x�,#li���vd��b�lL ,m�����v�BJ�M�+��Ъw��i-*u�sX 
�h.�0�X�lt�;%<��]<��N17�����Y�n͸��ﳐ��ұl#�,�7�}5i"��.X��[6
��|���"�����`�sy��3�@sA��L�YrW=[9���4��Y �5&7��Z��L��SծG�C2i���Hf��Db�<�"��|G^���:�,
�[w4��M�=��D|�=�X_W�4�*��� ������괫  �_,h6�8�x!a�C]�nC້Qj;"�Mi��d��6�E�k����4��w�=bs�`d��Q����̛�4I��������������A"'��Hhw"+��B��ɟC�3��% 1�軝 _֝aV����}�*�fL����N�U�X�"��;E4�f��r�Ɨ���eݯ�o=n=��LF�kyf�u�����O_QN$��� ���˔�-*?.ߛ�X�K(`��;N^ū2!NFʫV�0I,���wD�;�s=�$���'�j��^j��Xޞ��8�������h
�?�D�I���NG$٢�>�H���S:��P(�����T]�A��^"���1���|�2+q��| xߚh�4��vY�8�L����9H�vW�G&Ć�I¹J۰Z%1\�+͒�݆]F�c��_�OН�3|�&��;w�.Eeu9�}"��W�n6��?�''��ۡ5=��"������(��QuDx�������f0�������2��0�H�vTW�.:m�F�G�^C�OT�g�,%^�[������Տ߹��aC��Ky����6��Ww���Eּ�nv(�i���&��N���B\�s�;g*-��	��Mzi�Vg�/��b���y�r�Ά���>�C�x�h9�� w�P��"�GeS]^Ѽ�;]n��΍�(�'ѫQw�헖UG�ě��kD�������6sy|gn�1q�PԹ�ہ��2Dmg��P2l�**|��y�,tr����H��n�p��yq	� ��ڸ���dpϝ,0/�o��L.�����βP>��||�XQP	́���v���*�>�I$��C���w��`M�/F�\�&���Ó=��3��C�$�t8l�A~v@���e-9A�s3���s�L\�e
j���"A�i	�F9�R�VI�*4:.q� z�$�8:�'F�K�y��ɂ^%Y*�Ё�p��-�w4��"F'��?�R�:\2^DS�W�8���,�f�=?�-���n[ʑu�m7�Ur�B"�iŁ9���й�S�`�ζ1���i:�S��z��«��Dk� �輲O�H�*�\<jߧIbzت�aJm0�Y��ZS!R�lb�M�+��ujHH���
��?Rm�ی-��VX���H�c ��j/숽�a�r�!*b7�
��EJ�xU��%��Z���h3�^�o�0�=�1鷉l�ލ�  D]��7�I<�~�,�����噵 �oL���
�p��5�۰�q2��c�ġ/�?���P 6�2�='cMT�&���y��g(��.������
vJ���O�^���m`M��<�Ƀ� ek��l�{��»@i�ώ"e�
{p�=�X��Ѓ�b�����W��d;�`+ܞ۫h��(�C>|P�@دK�C��W�K�x1	2�65�������:�R&�H�����So)�A��"-qsɛ��3��`����@�;�<��Ln�c`AB\2+^�z&����Z��Tgh��v���ha���cs�Jc�о!W�m#Y��u*���케��d]݀wہ�\��b?�����뒵J��_�  'r1Qo�y��d�� �Cΰ�G_�`g�@zw�h�k8�>�y��EF_<b.� �#����u,,3�mmy�@욨�-2៴z����ٜ��>���CYL�#8����HF�_��R��Ɨ���zT��Z�p���TŻ�z�ꈆq7��b���1=UY����<�xXjΞ�-�d�!^d'��q�f!�
���̍Cn9��Dq�U��F[��}���_��P��,qMk��1u�sV-�Cĕ�Ԗ��Y-�á�xۍ
���Hq�\޵�Aڢ�Z&��W �&����!Y+����
�/�=ﶂ�7d�).��N�gK�Dm�J����d�{Cϓ6�ߪ����)+��ZB��e���9ҳǴg%�<y�|�KR2Id�EN�8=C3�{A�y��Y�L` �`b\g�Vb���w�ּEZ�O뢙�;=��t}N�������ƽќ��AK���
�(ڄ�.��_��
K����������^i֭���|��P_���k�2DI��O��?��%��έ0�
,qs�p�= Eۉle�A��!ڵ1�^�/�$��D��c���봥V���)�нB������΢���$l���Y�>�Z`�E������_�����
��n�P�pqi[���+NN���7wP��h2w��uh|�҃t�Hon��ASn9�4EJV�������}x�����d]5��.+� A��X���P��!������Т���bf��X�!�l1�X���O�m�j���C	[3�b)����B�����$�0�N�/��d�A$i����ѣ$O���8��s���w���ήؼ�.�%�np� r.�ڸ��Vg(Z	fŨc���8H��k�'�O3��G�O����+#ՠ8j:�ކe�\���穌�G��h��ɴl�Mt��h��&6�3�����ciꃏ�'H'q�gb9$A 7c%Wm, �C�Q�������ĺ������'o��D��U�9�X3{t�
��@(F�e>K��)����ֹ����ӁO2�mD$9wi#|!�UFّ��1�9N�����̼�R�Tza��,"�ղ4 e�g��Ә�q�2|	��g�H�d��{ �B���?$)D�BK�FƯH����x�og��m9*ޢN��gHx�oI9�5ӡ"�G�zPn�_�Q��K�݆�VЂ�N�iC��{!�Yw҅�+��� �G�'D�ID�i �t��:���H���U��Gz��D��c���xW��.q�L��D;�v�oa��S|�
bR�
s�����x���9 �s/��G<��8�x�V���߈�)[�L�]��2Ƌ������[Ok�Ҷ6)��Q��t�?��������;�3b�>�leF0�����׍����,����-W�5�S��kf�dR�Gޢ�T�J�i��������Plg���Zк8�� �R|E�? �Wzt�������
"�u����еiΕ�D�0��_�-DKV��.�νE3.F���J�E���1S�%�%��;A/e`��UEd8� AG��*��RBI���P�˥Y��`AyS�8��x�ɝ����ßH('��_�W[7!껅3�h	�S6�#�%֧�ha��y:R��<�����y�N+1��+N����;�/���/��
j|.M[�7ۖ��툹���A�`�G� �������6v�K����u�ErF��ð�:Ek�m4ވ�-+(F���$7��)f��6׍�O~>*v��?��4���y�E�}��#M�	�`�\5�rt��+�W�#
�,ʨ�[D����.��]}0�Kae�_|$H�ei���$����E��'�����*���p�ev��o�Gn�y����%~��Z�`�����,u8-��إ��3{�-z��\�h������G�ķ����#�/��U&�)��n󘮔�S��8�KOָ�[Ž-���Ez���fҶ��#�+~��#q�c��la%\��I'�!�`U�$�D_M�߻d*a�m!0>�QЁ��0�:A҉�Ȳ���{�nW��Z�
x���:H�����`|]�G�Mzk��Y�����Wj�w�?�d ��?��$���Q;´h�y��HO{,-<����a�2s����K��q�z+���
���e������÷{�b��n��f�B��	��'q�˖�&��d��%�&0��T;��d�6l�����%wx!�܆8��_�=�<�@4�o�nn8NCxG��8̩ܯXrz�^Rg2����f�+}�5��s��h*�Ծ.{��t}��_(Btk,�w�_���K���| M(�%�R��M�~�~��Z�Jn끾#�nz�	����<��j�̪邠&�,��BS���R����x���E�;޻� ���ƭ����F�!������"��,���ӗ]h����7����,`��I�)Z#_:��T*�fh�}���A�n%�b.�S�`�|�S�:�}i/���$7���'���7���V�-}��5H踙��!0�A��f̸72î|��~���G	����_z���׃���/�4^����ʽGP��R���U�ϸ��S�!4���9�l'����XXmB��L�b����Xc73�ÚΜ�C�B80���L_����dK�T'R�uhrGtWɓc�����

K���B����xf��QI�B�rn����"Cu�Z����	>�srZ���
�	�\b�rRx���Z�ë�mq�9��ޞ!�둞g	%B�
C\����o-�-P䖲=���YpC���$�NS�CM`ǹ��u?����Z� yWx%�W�o<�bgƽ�u��Io^���;1���x���cCh�TJ�#Q��6|��w���&Z�����,<�{������YMbXȤ'rL�w�dGH�f�kt����=���*a�`���n��d+�>+��V�fWK@��%��ʆ��т�2z��dF\ �Fu�~������?6@�֓��f ���C�i��˛y�L����� �K``]����`������ˋ0�l�#y̪��w���]���s3�މ����9�8�YsێwfV;��D�仗�ը�Ė�b5B����q�� K���i�ȕV���Xܗ?����4����#k��$\=o��
Z�V1���b/�jG� �cu:*7Y�=��p{(����rJ���A}�q7�����>"Q߰i�v\�Dx^`��n���I7T姇�~�>}����w��c�m-�$�;��7?z�
������fmB�� -c࿧��fÆ���Nf|9�lĹ���=X�"�4b"��
r�1��"��+��෰e���Ùg^�����X1v�WQ�m�^Q�.�b����Ñ4iG'���HG��[$���:�T,9��2�-�.<.�L�9�(ze��B���f}#��~'�K<�D?��*l+c��5)�.� Gm�!E�hf��1�tuX׼m)	�|�f��r�h���f�����M_�@���O�T����hy�V#e��t,�f���wV����q ~�o��}�wd�疏1�.�����<B`�$����=v�(K@�i�i�Uͨ�-��x&p~��E���.�72ȦN#Q��_���﹈��_�kѸ��p��A�1-�/���h���=����hi��g��7�����tu3r9P��v�cX܉��s�[��I��'ݯ*�;�%H�u���&�o��סm�,���\� �6�%.���=���|#���We-�b�J>�Y�7pؼJZAM�U�@���2�ob�m�
<Ar������0f�e�f	���+M��D�2�Q�H���T T�'?�:Q1/��-6=􌪡��n�b�}<э/q�ݐ�K-�K�m/+�ٽ�H~��I�S^~X�	�e�ScT�E�;$�%+��T>��8S^�Eq?�PԐBԊ�i�\؛�~
�]7kI�_�]�e�����۟L�:��`>s�{6j�>�`�|'�	bp3����(��Y��,ћ��9��]PG��y�V|32��J�҉���v�ȇ7H�r����G֊7��qD=�W�H//x��:�F�Ą��"��"P�h��!mP���<�*�c���\~�#>��J�W����(g;�'�'�]a�+��zŨ2C(��9@�$�5�q���$���A�uD	�|jN6ʔ�72�~�����ĽX<w�4�c�;��"����"��U�r� ?�l1����+�5�� �k����t+���M�z8�$�1�g���f�R֛��F+>�>[m5K=;Bg��= ��ؙ�-�*{\�s>Xn�F\#��_ ��(��}NUNn��s���'M*_k�`�	4Ƌ|�i�*��� E*1����W�M�Ӽ�ڠ���|�����X��)��U]*я$�}a��I}�xH="��%y�Bl0��$����׫Mݡc���F#��K��C��o�y�9������ӫY?I�kP�ܯ4���P�P�d�:!��0T˾op�Ͽ�;; p���~�%#®2Pz�l���WMa,�V��O?����<�������O��JK�-��RʵV��EH�"�m�)�R\L�;vc��`�	���	=��@ߝ�3XT�=��^�ԂQ����I�CI���s2�\�S��?�+�Uu�=�W�y�7
��Z�I�75������)J��2-X��)�ʎ5��Ty�`�d5؇+���%I��*�4VM��#�N\���C���bc$�=k�ĠL��T�#�j��+y�%�=x�V� ����Ov(��F����N�IH�q���O��V]�Q�_�u��F�a6%Q�+/��C����:��wq�ʙ���.�k������>A�B!9�i�)�#�L 4�Ւ�������PPr����]�R����"Kճf��+b�s���T�|g����˲���bXSڀ�VD�Q�!�a�aW�[fM��U�v�Ip�:�b7`�| Ԁ<�Y��)�s_�YVo��4hl�R$Ye�_����HE�B7�o�$����a�t���fB%iV�@�qf�̪�(N�����c��yQ6���[�_���
Y� �MK��z~�۵��0���x/
5Di��=���Tg����n{�C�xo ��rp&�zS�����f���,��� �MF6e&l*_W�ЬR�"�C��L���&��ӼTy#^�<���_ko��\��~׼�9�U����YD�>,�Ľ�5:�a��d��ʗ[�z�a�<��fP��s5��W��π�<���/A�s�G�l�G+����\��}�O�di��;��`b��(є�RN��W��Z!��k�v�v`�ݿ���=�X���3�a��e��ӃO�a������w���U���F¡>OH��HBFl˾aF�J-\�g�*W<�20�9���:�>�O��������B(>��R1�>��>t��4�](�������뽉�fNV��]LR(oT��7Np"�f��a��7�:z���u�l���M+�:X�#�Tp�2���|�oEy�O2�4�����o\n������\:I��X��pmg
�}����a
c�wcR�}7b}���\:v�]|�A�M�׉gm,��Z�&$J���j�c��h��
���wվvFT$�^�g�ڌh��gdJ��K�k���w>`fϺ2���u�� ������5�z��{�۸�_��E��p��[���pP��f��8w��i�Y� cuC_�dYv@�ó��Yyu��ޤ��
�o�I�q�y�zuA�g�ho��o��C�Q�_�YE���\��N!��}��?-��@HN���?@��d����h�\9��||!ٟz������w�<�5�7��`�k��.�7�E��LJQW\��ٞ��a�mU�E�l�P\����ǽf7�^�i�k�s�Y֢Δl��/��'y-�ю�,�_�n��牁.CS���3p�0S����`ɴ��7Y�ʲ�l����;��A��k �֯u-O�	�W��Q�*���S��ģ�W�����><qX���*���������])nC��G6J�ņm�ŭ���7ɀun֌ �*�ch�:UP���>����Il�l�C�d쾁���z�.��Y"��S�#ё�nS�����7�r��6�U��
2���k�`��$�~s7���eZ�%B;Z�mPuO�S��6}����"}\��%�(��q+]����c�8���z߄c|�?74�m9�=	(Vͭ��L`f��[_�d��p���{-��H+h�P��@r��;���7���*��q��p�p�m�in��������~!�<j�Z��X�����F��)���1\��x�FYӃ麘���%������.���y�����`����< SM$���+2����9 
D�`�)a�1�6���ȴ6�� ���˨�8��2��!�@WË�HG�V/f �4�/��RP��`i�v�	��'��v�#I������Q+,�J�դ�p�mkT�[�����C#g���mp��h�����4ϲ��J�#R�oK�yh��k6�[�A��?5;�'_��=�d�}Of��C��JƲ�ͫ��^R!�	�0MPa�F�In:byu����6�f0Ia�N��df��[�.���O��8�����k��Lm��p���]����yGe!n�ˡ�h]�Q���k�D��D���kK��Y����1���"wzĐ����,�&����!EǮJ�q4��˴�ޠ@$�]O���iu?z�&����H�:����p--)Ϳ�Jjy�p��@���K��]�*n�A|J�\�:@�����X%��;���1z3�:n����r[��I���3��>��1_�ˮ:�H2Yk:䗲�d\�Î�9Ƭ^���\�/�N���>�`r+��C0�#�)���.6���a⨓����p����s�F(�cn�.�"�pb(1�l�缋?��~���b=�V�D��� s�֞�i'��c�W���P�7!���M�+R��ȝ��~^�A�&sŌ��=!"�V}�H�v[�X	���qZ��G	j=��k9鬒��"�K*���й�5��p��a�V�Ї+B�&14EE��$�&F�xҵʊ�%w-����*���2�~4U5���.&�h2e�|���8:�p�?�%��Xm�a�j��̰ļT>�X�Gg�m��*&�~qW�y]��i�(��l����q�bA��ɮ���5{��U���I�!љ����,\��I��E_W0H�����������Bh�k�8h�ղ��)ב���&C��d!�&��uўX.{bÇQqk�_�F�)P�b�z�Ajx�t<^�CX��f��6|�Fg-�6�",s�F���fM\8�։o��O�&��>����;�2��N�t	�``S�.8e��%@���&g*��~|9i���}1d8l�C\\e��1��k�ʧ�9�g��-��|�s־t�k!Zc,�m~�}���@�g�}����ƚ�%Q>��{�H��%�	�g��g���w���v��o�AN���q4�ܓwo�{���SK ��`9�98��7;k�C��f�Ѱe��FF�t�2�h1� l߼ܙn�Su�c���5R��`B{�4���-�xl業�;�)�A�~D�kVb��"w� �-�1����~aV:o6�ٶ���h���2��Fĉ96e�+eX��vS�/����W��햞�g�la�2�6�Aq]?����RZ2�(���h��}��Il?��2���(^�Q�����B�|�Wk�
^.��$Evq�����NZ�����C>Sva�Π�́*,��&L���%#�G|M���]�!����7�K7ӟ��ӥ@�}/���DK8`#E^�:Ptv���WQ+V`�`(�~w�ߒ	߃�K�=v6|@VO�����>�K��-�Q���^�w�}�txk~0�4�pl�Q}(�-T�c����n�����b��{���/7	 6�5{�͍1t�)CM��G�kU��،�䕼!�����H��.���G���A�]u0��>��ms���[@}A@�����q�k&�eZ0��?�w俫m*��,`G�P�]��'�,m!�xx��o���y��pl&������N슈8��{�P�0���B*B���a'e�"�R;��<r����fj�����t�Ĺ�o �t���5����H^�����[��Bx�*�k��TF����՝!74|Hq}Y�L�<4Q����p��O��1�
�0i��r��Oم-�:���|��`�������r1=��=�.G���6Y�{���i����FP��Jހ�l���ѐ���@ 1��Z`ڒ�d�]vǊ�U��kV��UOM����+����0�)�Lk��g<Rݞx��e�ѣ09�1��$��/�r�\U�з9�E_`��S��K����Ci)���#tɴqE��N�\����!�D�Z~ɛ(�6�-�;�lU�mE��|>1�M!�kR��Ub.�����6Q�v�y��H-�?x���a�|X�)�Xݾ���h)���>��g+�9��[��'G��}:�P�5�l���x>-D�We��#�;�".�Mo�_�Q�@7�a]Z�M��k&�B��("8[j��Ѵ�H��oО�����w%�U6s(�����Uן�Z6=̄�{*.�K=,��8S O��χ�,>՚E��:n��)]��*���N	w�w�!�=��Z1Qs�Ke� 3�8�t��d����04ZΥK����p-Q�m5���F�hq§HWB���ʶ9K�,Iݛ���n++���(4=�'��j�-�f���P
�20Dͻ��H�A����|@B,�t���9��uo��yJ��[�
Pt��U�(�����dbI��|��%X ���ޤf�7󫏋��
ԓ�"/�A>�%��3J)��uV:�h_��u�H���h�G$y>�����bGo�N�C��@�C���]	xK�O�_�)�0�g]�{B��/�w���w�Lb,�B�3�=+�s��mWr�"z�N�u��[�t˵T&������<'G��^OM}��(�RZ���v�*;�-c[��Q�'9�?`�z�st��u�n��Eh�S:[�)�ZS�+��+8 ����'�-����
.[iP��	*��a�7$����&nX���%!٭*�[�#_���j�x��a��E�
�Tx�����[�*������[���"��� � ��d��6�	��F������g�Z#3A��<��r_����Y���*'�K���94Pdz�.��z�W�i��zRV��P/�}�mg�)X��J�1BjxZ� ��x�L���A%i=�v3�"�.�2$�Dd��/�|޸�ev��UW���M켰.3(��k�F:�����-�|�|�Pk�;D��ʴ~�#����Ih�~߰-�ps�6>י��~��qqT-���Tx�#+�TS眙"E��(��!�O}��^�VlN۩������@�'�nŸj�Ŗ�=�S�U[x� 1;$2$�W8�q�����K�����E��?��J�a�E�O���8�O�!~j\�Xg2�o� �
�c�%�/�N���{7��R�fa옣o��5��r�ҹ�����֖�A��Rf�Qs��5j^�z��K[[:�e�>w�٬:���Q)
	@9���BZ�k9����i���0��wᐛ��c��4�zY>��k��K_�8���9"�^n�v=��r f�u�n��;�aR�0��!��^�)u_����9���4{�t�7ֳl�;Ȟ+�r��� ���h�K�]|Q����������tD��;�E��21�� �����rj�VC������O�ٖbC�Ɋ��B,���g�in���(0�5��c#�k��'3E��F8+-j戳k�����d�0��ߑ�}?|=���S�I1� ��*���A$c�܇�?�I
��eF6u���V�gyV���h�x�	���z
b��
Lڟ��
�P(�q�X �,�lz=�gm��r�,H	���j$K-��������>�3%�9���bGV��}k	����kk���/O�E�V{L�M66(�!�&�g��7ԁhR;��֖��ѽ*�����\:��OZ-B�"\R�܍o�y��u0h�@�t�p-|���U$>u���|���X���Kd���R;�d����֎T�&o��G��} ����whm1yPMO����/Q ������]����'86���)�T05Z��5O$'�-����A�(�w�N�t�gu�
��r����2�:�:�Sf��ȡ�����4K���XY��
�ţxi��R��;x�8�����5� I|��I"��1��/�����I����Jl�8�e��o���{=�>W$��g���o��/d�G���j8r���[C8=
��1^V��'=n��C1����.�$۬��f,3J�[ū���둊O=�����Ad��;&�%����(�%S�@�D�l4���l�ǆ�3и��J����C&G���μw;��	f��+���^�}�{��j�o]ޙn�Q�?Qj'��,("���C�O�	�v��h�cU+J�u��΁G�L�nո���k�{		�T8��kbN[@�)���2�R6S���Ӄ/f�����Es�+��Lyxo�8FԌ���|�����?���RO Tߠyk>���5�V� �g�̜5�FV�%������L#��m��W��K'�Ν8]G��I���.��i��;���U�.<-�Yb(�����^�|��'��=�َd<�aG|pX�Qvd �,�yޑ�>E�)�i�F�=�/�Te�"b��d>#�̥�y<uoN���`���]ĂPV[V�fsQPf���nLϬR0og�Xٌ��,��w���v�� �%s	�qF���b��?�}�Ac�R�����E���/C������}��e4rE�x���:(<�]���A/g�>N�O}ڶ3k�/�w\53 �|l�h��v���`]I<K܏^7�r��N}�>��Ϻ�e�XB)�C�u�q�܄��z�\%n��sƗ�֡�k= �|>bTܙ3�؞��P$��x�{�yu��O�?���]�RS������� oݪ�/lP��� V�IzO�*�['���H+�MR#U����o���ύƪ�P�J�kY�	3���c�f���Af=Ъ�,@����/���ǣ
�D��!ؐts>���g��~c�'��$A��#㭔@���S��P:�$�]�w$���ݫ�؝�TӺ\�+ z��8���?�����N�$A�Һ�����%���R�f+jz2?Ӷ��{��όз�N�|�h�&��pl0���]��x6���l�s��~�X�.t�(e�g�k����/�|���oC-�e���TV6M�t����yU���QR��>	����zG���C?���e��G���9�DT{Y�&	V4m��`�ش�������!�`���ci
-lT�Z��$�@�pIv	qU�� ��^��2"S^$��e���QFkԓ�Y
��� ��t�#��,cCn�yo�`�껇�T���Q�gA����V%B����;���nD9:ڹ��xa d�%�-����x�h���l���qLϊ���4Oz�v�.%w�1m��}3h��8hr2#�|=�]��8�ŗ�6:���
�ο��n�/�b�c-@�������B��<�Eg̱��n" �+���t}��&0������z�JUt>&�Y�>S�b��w[�E�yaA�
��'+�	C�E�e�:�遱c6�>�Sd/Ӛa�����1	6Y��͓=$����W����)����?	�e`�ˮ��JU!<���ڸ�9/#�c}R����e�r%�ò��8DE3�u�`���}?v; H�/<�'�3��Q&�4&F=Ԃ����K���ŒxA�b$��_��~�����Et�-m��w��ȓ���է���ִ/�[$Lܨ� �|���82u�W,�}��=�w���Ŧ^���٨ʐb6���4�{5�5R�u�X(�J����b/���($k�������S2`?��y�����u=ژg[4O����~�r����fdP��8E�4���5�]�����'��W�I3ҋG� Γ�b��vZ�;H��Y*��U`���D�|���Hq����(E��C=ʧA���.�Ș"�O�8爝R�Eew����*�\�OuW����e�B"Z.S��}����/�QNY��J��]�{�}��`mV��y�H�����^�O4=a�(��������>�ӣ����61�)����+��0���or��z���|h/��a�j�P����P�>?�A������I�!І���7E�ɮ--c��w,R9 �h������0Ð���s���_�=I�<X;��>�*�����m����I�t�����(БŒ����.�B�V�����p�e*�&���Q�.�hpu_Y]G���i�1|a(��T�"�ěA;�i��EA��u���cJ��(ρ,`��}������h"[��/�y����R��_�4��$7��0r��ܨ�7ܽ	l��Ȯ{�}k�A@�"!ӽ�l*2�^-���20�l-?���d�l}�X�a�"�����	|2*-~잭)�ML*��i@����_y�S�P;h�/��1I���͔cg�a��,\��	��I�y$R[��Z��o�!ߙ��EZj	��`S_?j��F�:�{҆��+��CZo�ho���}����wҤ�wQ��v��h�Z}��> "�	�g"�6s6�o�uц���|G��B�Yz��i�A�I�<�v�fIW�`V0"�M;l��m�^r����F3̫g�  :�i����=�ν'E��# ����Ԏ���-�� � :��A�y�~���S�.��R�u "z������GqUJ���hB	�T���8���EY��eͤ$�.졊Y]�b& =�?v�7�(%�t�T�V�%�W�Ԅ䜦YD������9p�V�w*�
����f>׳Xњ%Q6�g%i�C��c��q�`|��;���Toa$ip��dP�m�Z=�F��U",N"��y�k�,�AE����gx�k�RP�ٍ2�'p"g�u{�P���k3��&2���Ɏ.�N}DO�'Qt�u��E��k��B���7���y�+�C�ABB��۴ƅ�Bgm�-�]�R_���)�,����`�D�Q�b� P��t̨���ޖ=V�NK��zW�k�w^I'.�r0YL�������ҿ8W�%�D�r��/���t��Tu��(���vc;�y|��P;�1f/z����w�V)�?��Z#�@�llQ�-m� �����(71��?	�AK�o7.\�y�Ȟ�[�f ���$�n�[���&�O�@n΂�h�-�l��WF��1�D��<]�H5�Jrg�\Q��X�0���|��n�������������S��QR!w�{En�YpՍ]�3ǚ2^�s���)���ޛ~�x$�]oCZ�:��t�I���3L�Wg�_|�0c��A��!6�Ð����
�{�[����_�^T�����XsoB��iR*���M~�9��ظ���t\����TG��
��� ha,	9mׂ�k��P@�I?�Ҵ�`b��ҽ����h�}��9%��T���`�پ"�ŗ������}{8L;��k3�^��V�)�����tGF���X��,7���R��XsZCfB ���N�W�&���őrR��,�_� ��c^QDR�Q��J���"�D�<�]�0	4s"s�!+fWd�!%2�^X�q�lq,�Q��7<o�\����t��=?�������C�Ƙ� �A�&��{Q�#��S��`o��9�qǗi�,�Ƽv�cW���ǚiPE^�����K���.$_1Â�ɿӂ0JE�PZD�����X�!J�0TI_hG��.�d�_� ���܀������_Q��Juh�Ä$�I�R�u2m�(�1�*�PePa1��п~��c�L���ޤ����Z}���4~���E�s8/�{�=�-�����gJub��kgS�u�s(��l�a"�8�D�O�N'M9�~	2,9���������f�YY�X�0�~��SMc2悀%z�gjK��ǹ�;W����I��:�J�"Mu�6�iS���t��T�q�g,E�{~"�,�?��\ ݚ��r�~�z� ���`��pBV������l�}�
�~E�JXmn��h5Q���v%�=}?M��E-ls{t��S!hJ,e�\r5B��~s��<�o�Xw�\���c?EJ�*����t 69��ӌ[�а\-ƌ�^���J��~p�=��d�n�QǠ�/�vm�J�e��
<�B
q�u�b�gz"r,�¿VOlHI�e�jq�N��B�tL� g�#�0KD��+<����rN-�za-*Ժ�.b+��R>UVI5�GP�y۷�{��7�?7�Wn�_t�?Q�|�-1�$Z�# �M(w����$�\]ɩ�XP��L���DI�P�SpyJ��SRvW���;*���CiO��A&�yj����� ���Ղ���>��6uC��v>��c�)Æ�����l�:�I��Ca�F���5+��rR�޶��O�����>�~M��f��Z3%CV��'���-:̂�����޲�q��7=C'��'i:լ�0�H��)AA9���C��g���@0�G���hB�I_n����[e�1�wWzme���˂��Lh��&���� ��g?G�P��3tE�գ����_�Vg�6��;�)�Q!������ �XZ�� �Tڏ������	����ae�$��RF*��zcԷwQ.lh@	����	r��D�z����w๙�I���5���H�#�yx�Y��s�^_ީ�n���|�ޕ��&4 t���	�q��C���5���eB-F�;���2=��O޽�&���_w@Ǭ=�y�𻢳�� ���0�j}��'˚��8�"7yɸI(RQX)q	�-p�l���$�&�un�����u����X��Hn:7fs.>�?+u���g�)�G:R2�0g����݅1�(�	�*�z��%�Ԣ���~�(�n9:�F�?������wu[��5��u\O��&��)����2҈&��KQ�/v�iSgm~*�J�C#ԝX*}	�-~f�,�*81$�?��g�vQ��l=3ܽcCY(	�{�'��ufuN'2�2<N�\�j\4;����]���;�p	Ŝa�w��;���JN/
GJk�Xy�qI&��� w�V��0}#3W]�a�C<�r���X���K��m���[�t�B�i ��A�(�m��V1e���5%Y��	������~��|����d�!�1x��M�A �s~C��Z�Eo ��3�]�Go��ѳkR�"cRɽ�E���Z��-o�E�`�|q�߿�z��&��R��&����7�C�AP7�R� U��T�����iR���P:e����Pؖ�t~�Ɠ̐�E������>]�W�A���nU�*U�]�&�?�����κVM��:�͹��_i��\k���=l0�Ͼ8��*��'���6���A��z<�ݚ��D��`��KO)��_ю��"����]�8}�h�@;���G���V�g+$�SR�P�Y�q���t�'�ͧÁ����,c1hn�2 ��db
�9�������q�3S� �������`
Ȥ����k�j��=�D>������^���Ҁ}8�TFP�v�1��q�W
Gnj��i$��b�ȱX�X���2H�,�
� bۢMp1�q�����Sؠ�j��_��Qߴ܏�K������f�|ً�r`|NagE�p������3ͩ��w<�	�"�E�r*���Lf�T��7��%��pk1^���Y��:�����T+\��5-v�`�x��t"��M:�W��s�KR�����pʐR�#�|n?��N5�����2i�R^#�f�	Ҧ b1��K!܀T�q�ЦX�K�k�d�L�4�@��nf����q*�)��bԙ=d�P	@������5�8�cɓ����C��Lg�Gg�c��<�%>�y�%�D3���Y��{-�nޟ��p�n>��d_���k����i�[���*����������k�*6���2t!t�H{�[
ᄛ87Bik&3!/Q��-�N/�6�L�Z7�9��@z�XQ�P���P�d��;ۈՒ ����%�)sח!����+����oǄ�VM��T�eC���ik4\$����X�W®?1I0r�=�Y����&�x�ے�V��{��p�E<�F���B�+&�@��],��� ��9=� T�-֝�ۃ��Sm[#A&�����%��õ�C˒�IP"������w�ߎb)�8�-�^]/4��n�*�)�r;	�F1ʜ��0̈9�Y!��{s��ɩ�1c��S	Ҿ�n|2m�Kk�]�|�&���FL@�H�Z\Q�u���hn����Lyh����LKyX��BcK��P���X�Qm".��/��-��;��/ʈPm��'�9��3�YD����j�,�<�d���;'�����K &��r���H�G��a֭��$��oݘR�OdO��U+��7���ygd��7� �����Y7�RZ��D�5��maJ��F�$`q�t���a�EE9G�]KC�S�~�� ��>��>iZ�9C�������Hb�3����-��h�9���
3"-S��M���,VIM�iˌ]�m;��=��od+��h�S����R)���V�C��."�o\��L��Zy}Z6}%�:���#�;^h�j���"���	rg�B.�vt� [�r��u��p���<�q����X`���_y���l񡠶ӑ�Gw�^k3.�.���j�ԅ�����n\H�;�eo�k>�T��ո=ϧ�p�,I �5��,�|�����ҟХ��Ǻ����\�2W���5��=���O�ʽ�pV0�D�?���t1�	�˩�Q��2�<�m��ߝ$=�ڑb�0�xV��3�0�m:�g^�SK(趕^y�D�%��>A��]i���6����=��k�P����I�nĭR7N���/��^dp��f�����Ep��/�@��]�s�p��!��{Q�>�9��1[�������,���D��!��jZ��w���1u)XD�kX��W���Y����h[�^A����~�RA~KńZ��xg,]�[o�o�<*"&��7qT��;��\g��S��4$��_[H:�9��t���
�Q9���H�g�����@0Y��E#s�w)�XF��R1��kW���E1�r�1�1|��o�⧊���ǝ@��ꓷ͑� m=W�$g"g
E�} /{���B	��j�3��O���gx�5��4�b-kc�=X���m��i��9�>[���t6��_g���|�$	tF���eOS�^Q"�+Gym� �$"�O]�L�^�F;p؂�g͐��N�zb"�zS��FBq��*\}-/K���i*�Zk4\�(�n��֘��H�����@r���uO�,��/��<d���D@��y3���N�ᡝ
P�[��险H�9c@�;��@���_'y�34��:���:�Z�J�\]���c��e7�F�69�����r���l��Y^�4B1/��?��fB���G��V@�U��#u Ę��65"S��_���,��a@󵩌�2� �|�߱C-��t��I���� a��"���`y�}�hZ0Y��Z������m4ޞv�w������Əh��f�L�����3�څr�}C�/��f~�/
sB��0�R�[�q,�2}��~�(֯�u�e�����p�c9�%���*��K�*~�]Ȣ5
:��;��xn���M˕e���9u9^}2����7�iS	si���˚[�m�D/���:��Nj��Ƞ��Kt&���*cb�a�L`[�@��u��B�����)6�נ�}�:shQ�+ݖ5\ �۩���TZ���_��*��$)���Ӷ������_��V>Q6��{�i6k꧊S{w0������h�p��|<��I!;ps�(L>�I��H�`s�������u$�%&;������a�K/�i�T1]�x�y���Z	�;��%mON�Υl�>��!(}4���h`S��|�A�0��W3�ZW~��i��9>�W�8u�ٞ�<N�`�rR�V�U�|�U
+W/ �Vq������j ����0LGF0~�X���`��Q:pm,J�ô�8� ǥ��Lj_w���n����z�MT�<
�m]�[����ЍOG�r�
��N�b�#!��!`�N�꨺�Іڌn�Jn���Yz�V��w7�����uKұ��*@*�o�>{��4	;�0�{�J��F6�^�U�Hg	�.(T��z������pж�N���i���`[�m: {�	�U��6vs�Q��}'�����b>J��0��iz����ߟ��Y�gl��]�ݏ�.t�.O|z6D1����JD�:Ҳ����ja��1�)�'R����V��x{������� M:p�O����')\#߅d��|�3��9���Ğ�i8m�V,�&�L�8��ݝ�ca�~���3��z(_�o#0Zj���~�;��T��Zn��ݟ�u��SyJ^G,���%כ�1S�n.�{|�|��x�3N�)=�),�n�!F�M�\���\E��|v�*�-�5�cv�d�mJtmT-}�L\���EYc�M�?����������0|9�V�ǃ�96���-�х�$�����B&�H9�d�:nT�%�gl^*	�%W��"��-��7����-��`�*�&Z]�������8�(qQ4�h��mdM��B�[�J��ȳ�a�H~�������A�����x��e�ċ8ѣը�_V3�I����L"�@�{���)��p�}v�4W�����i�D=ҋl�KY�s�돞����P�#��Y�K��p�P���wP����"-�I�m'�����akQY�VW=���wfSTTu����Q+"X�Z	�4����Ѧ��y�͞���t_�H�y�=��ٓSGj�"�k����o�i��bz�x� k{�G���}=N �!E��>J]�� 6r���(f��H'9�����7;k���]���y�ȃ�����_�K��PQ8�	k�F�y�+���T��3�fVx���3<z|�DtX#�Q�Y�wݚ����Z���v����N�q�Ɨ�3�V��P�/�=!��{EE��ٍ�sdm�?�Nnt8F��)�ET�S����-1�/p
�H@;`u3,�ʢ�b(�b>P(�h�	���SB�"�efa1�F� }�wv9�k�����P߹���߷�D*���h.� -���0�D��B8�:��W;�J�XnC���)�}&�m��X?2�w��CP�?���O|�Q��� ~��8�/������Sf.V�&Ĝ�FoD�*��E��4]L�``�8I���B+�֍hv���?�C�Ϸ�(��U��M](�0x�'�ll�S�f�6)<��?�K	u��*���s����M�o�5UV�H�M��c�E�����S��͓�녨�A�/�����,�ffJ^��������k�D�ϼz ��+'<�dnl����`慟gb=�ȇj�W�p���'��4�,�$�oRk�?�I����aa��{4r��OlN�Wu��&��S��\:���Дh�}���ȣp��>�O���6�w-���MiH6�s��~�-�14�@���:/8{�Ք��*㶹g 1*ё4��$��(�ƻ��a�u7Q�~h�y�p�)��H��A���&�*�"����=�'��������v�j5]D���~��<K���\E�b�MAa����Yލ͉*���Mڦ@�Z|о�L< O�U�6g1�+�Y-6��4J
-���ݜc�p���L:NN�����F�抃�x����\tb�!��-�q�y9�HI�o���o�_,1�� yw��1/j�������!�AX蒈(\�s�A~�%�/��2D�GvX���Uh9%���E�pv�x|ѻ�al�;�����(��G���&�;`v�@[���ٸ���qhKh�/t0�/}�L8�H)�%�v���d�S�DT��bMG�3�-"ґ����1)p�5��ӷ	t�VS����XB3'νg�*��(�=��#X��z��ƩH|�a��4E���@�hF,hD�@�7������;�,���)/X=-��2}� !�;`�������̀ԅ4�IrXVT�b7G�ۤ}~�V��������0���L�� ����(�sz��<)5�@o'�F�vP"&�Q-�|Z���
�֜]�F���B��+MJ��'K���"h���K(�u��R���@�D]_�ﺓ���c=˖q��� �Go�u!�.��)6f��a*5�װ�bkө�K�ڮ�
�n����
?k�����4����ƅ�y\�T��Ͼe���O7C>OHQ9ؠ�|!ҷ�kO���R~�9�Q>2����/�^�0��Z��~�m�kh}	Q���F��i�?��߸#���'�O�Em��|����҄D�V\`4�|F ���d�xg+MY�[�V̂:�!�'�S���� �����"[�Lq�55�q���'l������5�P�+�G�H��G���LTx�ws��E.0��%�A��x�(�=���;l	"�B-wv���u�..]�oo�g+��lw����3�e|}�ކ(�p�V�ni�5���vj=ZN!����崯0,s�~)���"�\�}�Ч���+��S,ꁩ�gC��/P�@b�2�V�ޥ�����N��x��,��Ziu��cӀ<)y�.:�f��l��ܷ��W-
Wh�]��X��� X(�0MG@�+�;�3O�Ȁ0g@	�X��T�J��A���D��y-�RG!<h��:I��3�vt#7���׬w��^����`��t�� q6(��!��e��I,;L?��a�{�X�IE~�9_��@��=�eV��c)B�ˌ�ă]���t�U��?�y�vSk+b�Y�q%�C?���x{�w3Z���'G���|a��:��s:���o!*��:���O�t���H�$t�X��gٕ�
��2�!�SI�6Сp?��29eߡ�^��}���'VU����r���h�Mh�1>Dp=�QN�
[��:E��#w��ۑQBL�l[�2�Ɓ������V̆�ӄpe�ao��~���=�+��XZ��'?ӎ��&�ߤ˰����{O�rٞ����`�3ϻ}r����������0�F�$�`[ł�/�z t�N�J���g���7☠�>-MAj��O�SN�����4Y���T�8P5+lӚ�����������Ó�6�^��JG�p���P�+c���d=yGG�A��d���9�f:���m]8�g��ܜ�����BK�_�,�3B�4�hN�m.���f�/"�+m��;Ģ�X��	����<5��]Ծ����'b7.�"�����d������M�O��|h�����4D�`���
Am>֋�Ss.Kt{��_RU��F}��۵U��z� 0��̶�����ݝd�Ә�т���ܠc�����?����0+;�ke6�8,5�,�M/7�9�� 29; ���ZZԮW�1Bk���3C ����U�{��BWX����>=/�b%���B=�!W�*�v@&��׍���K�%�UȜxc��S�&�g[R��Β�f�@�i~&��>#�Cj)�2z��r���x$�T�wD�F�w�F������~���WN���f[�j��S��	X q'IҸ����<�c<C�%xdL�6\9$�I�b�ËKD8S}�sn0e��q�98�gY6��m��z�m��jæ�Aۖa�o�pv�WHK��)���䤔Rx��)�Ҭ�����BhNĆ�?�W-wt�C��N�殂��uFND`�sa���b��<�y u�:���T�-�q^R�p�l]�ņ(z�攅`�V�y�,��t$�e����ŚM������O�OG��}�˄�j���t�kk�n�˟�Q� B�{�3�VAd
q~,�Ҙ�_�������R����@��=A�J}@kf��Q-1m��r]��r ��0���"a�G��Δ]D�:���^������._�"Zj5A�%�r��� R
 };����(��L��R�]��g�j�M���a�d�8H�9:%PxS9!o+�*)�����Ǎ)&��܏İd_S��XN��\g�FK�@x�l!��UJ�M�����2o<S�bO$�kH�u����aS�"���Q8&��[*��f����p�Q����U�shai�FD�le�� #��_��(��>X�XY�v�_MR�܈?�������?��م�s�ZW",H?N����H�� �@�k�X�FQ����KK�l��vA�\o�Z��&~E125���kv�����U�������7����D|���!k���|��i��g��>Je�K{!��_����b_��K�@Q#� ��#��x����<���0�>���U��{��h�Tq�+t.��L�{c�CZ��8.��FO��\�$]���<r�U����f���Uק�] ��"WO-N�/j���8c�gtW�m���A������������6eI0^]s�����FȦJhyM���JFV?-&V�.��eJ\�X��s�G�}�_�'
�o0Co���.����_
]��V�ت�XUs��Q%l�AZ�\$v�=T���F`=�Aj{-󸃽��uCw���l�Y{��#Kx|��NW�&��pL%�����u���%=!��%<AG�F����j��Q�{BژU����p���"B�X��.�˨X##���!��4e��6��7������_��,��D��&~e��,I��z�l�%���c	χ� �nB�I��P\��*��X�Y���i�b�b۔��U�m�'�I����tK�m/��[ր� ���e�5�t�8�f�{5��T�ޠk�S(8�	0An���j#�Y���j$��y�DT�|�fJ�{e2k�����b��G�:9��N����C@�W�@�����j՞��#V}��� ��>A>�L��������8l��Z_�LE���j(�2�^~IeǨ̈́�H�"&�2��v��#��0׬�D!�&==�O|U�o�;�sl�?7b�p�o�ݦ�����xv�$�emCk��h/�0/�G�P���9h@���X Y������$��t��i���r�T���"weȦHO2��!Ĵ��{ra���'��-�y�"��k���I��(��cH���8�A�����Jb�E���*6�b~�?6�ĝcf�����]g)&1OEu�^�{E�T�j}B���[U:1��T��1�����׺����x2;�z�$͛AU��?~�O���<r���I�,o�P�2������ʕ�վl��O�qi����ʔ�4�!+ ���j���&�S�q������������P��6t#��\����8��Ӑ��;��H*���]M�/r;o�0w��3��y?Z"����I+�
�5�n��%�M&?�@^I�{��TCƌ�b\x��6	�T?Ԕ�Eu绻Qv%i3�Ỳ"��^�P�m-a�M�{
-�b���Gp���a_$	= ��w�	����i��Ad�4��
d���
���ˠ�/3/���d�C(a/��趺�+�;�T���&���ґA�u��~v�w "��f��2Im2*/�;��ȩ��5����I\��Ձ����f����g�$�>��u�^�4���D)�1�1��5Mu:)�^�����Q��k��)=���^���������%�ދ �����q��c�r�`�5�񪌺�
��� �B�n*$���]7- ����n�P�d�PԛWSgY	��ԂNz��~�	�2��yX�O]�s{��"R/��ˍ9���5��o���j�5�r>z�@	#Wid>ost��ؠ4k�ц�+�6/ݺ)�_Ow����C�j[�h��i�	DU�unL &�������a�NE�xg���@�4��pafm>����O��T���(�6��AT���`��RxN7q��d�9^����}ZBXyf�?Dwi��6tu�s�l-�4:GJ<�i�����c~TWAZ/�-c�-Pɳ�m �Ź��yE���A�Ek�GZ��R��Tp9�KVe]������e�Ǣ��'ͦ�X�26�G�t5N���O���^8�#Un�E/�b�d}1	�(���q�CS�a@�IgsE�G�cJeo�W����]�����F�2v�����q�>��#�DI�#z�c��EN@7��@Ko�ot銞gd�?Wy&��I�T$.dZ����?%�l7Ȇ5���i�����֎�l}�Pۊ~cR1"=�w郯��^�mA��C�}�N�VM�&Bia����</e�f�CT	�`h��/��E¤2�[P�s)��X�'��B�&��X��Ńr��Z�Y	�r�B(�,����j�[P�#1�Ӏ:�/W�^e���b^_����R6�c�.Up3�È1YS#� f�9����_�">��pd��f��;X(/z��,�m��]�=��Ѩ!�2L�"MD��S8_�b��[���i��8e����p���Z��:�xdZuI��q9S��z��������L��'��I�B;�$󕰕���[6�eg-�x���y�[(~�G�9�!>���Uꔩqk�[�1q�e�74ҿ(��ۆP��1q�,�햋s��O����6��^�C���!l�>��� ���.)P�=�q��O�ކ��%�p>���-�9��܆�p����8�������:�&�ț}U{H��AH���僩=�r��FT ���2��A �FX<ke��!� ]TrN���BLJ��<�@�����m�o��E����Fk��1��7+�q���
E,���8� 6��r�))��A�9R�pl�Ut9����=,*�W�#"��F6��ʪ9��g��ǣ�Ak���ɘL���f��>p�_%�lʫfU��k�^�������[�Y�'ϳ�Y��>�T`���`�#�Yz�]F��1����)�ї*��~]��d�%sU���l���f8al��J���h�pF�;h���W�?V�Y+��G��h�fZ�O{�n�ұc6�� Gk�^z���dR��hf������L�:n[8��L){��W���E�XZ�2A쮴�d�G�,L���k��|"��qZ_��	���; @�BJ���ƪ���T��o�.v���]�i$c���X��mp���@� ��f�}@���OV(=Z4���\�~��y���(�E����=�a�Ž2���t^]���G��F,�D�sD�f���F�K0�Ҭ��oM7$��ݫ7���� �2FSO��k��/�_W���0d/l)fhVW�(l�?[m�ã$�1�Z�*���PV��$]�j�7;��{*�=�=2����~�Q	�i�%�z��ڏhG�����
,
�������<!R��W��L_Es5_S�zO[y��D�ړI�@R�%@^^�`��}��]X1�햲Rr�It
�\A�n��`z�	'�\ƌQ�?}��-���3?���hR-:��Ŕ��z���VaSz%w~�Rd�|@�������I�F�n�-cm�ʕiF������ѹ�瑙2-U��e����8��5J`���� �s�_��Y�y��U9�Y!���7�1�F�Xm���f���&&=�M�zσ*�%��̔[MR�O=����V)a�-�(��Qu[�3ת��fb��j�	^�9�Xh[y*��sߏ踂?lǣ�iJ�0�s ���x���ғNl@�\�dDJ�^����IU�1����-��+���//. 5�a+d�e���2���Ky�MV|�F�6	bԻ�I3�i�}m�Ȳ҈q�Ƴ�[(\��Zu⇼���u3�/�
JV�q�*b�1����?�����
7��.��P09X�E(=�1��~ӵ��{�i��e���T�FI�.�dǯ_�)�Z䨔!���Qv�_�c�s �0��h�dk��v��;�3��-�S�P�N����Ar|�����OTV��G�9�b�{|GŚ�	"U��[L��}.� �E�M�X]U�ZCl�	�SX<WK=o����jN\|g�3��۳~zv>"����U?����x�֋�� ���W0���C'������l�B�!V�Ǩ�J l�Q�������BΙ��i�rI����N�%=���ô�ߨ{nr�e\���F��N������3YM?'#�}��TD���g�<b�L;��'`Wv�e�D�/�x�T�8��Q'�lB���l�t�{-P����D a���o�ď�5�s���6%��ϕO5�s�	7�Rd��r��#u��G>����t�"�<��2Yd���mHФ��7^��ؑ�O`+VSA��o��S��X=�E�������7��ks�Yh�>upj�)rA��Dr��[�I�8��^��@��T"5ayM���[��D��^�d�/$W��r���}���L[ީrC�	� �-�a�n�AE�+���������-�Nn$�j��dEDev����S�o�R�����ڧd�S�4jE��-����i�>���)J�~I��(L&�4��/��W��iQ]IƉ]�p��8��Jr�C�į���	a��n�_6j/�*	����ڙ��"K���U'*���Bh�[�{d�r�^������~�k�Oi7�L#��7�F�`�Ц��#`�M�NG����GF�e_W���g;d	�p���kc�2<q4��"HlI��F���/����#��(��g�2�� �
��y��7�Z,�������`�u@��A�*���1j���>��lt��6�nc��7˕R�����]�_�i�?ơ?ٛm�2_;���2��5N��ي�.����N�\���b�<�@���X�h�_��هD�s�[�8���W��U��IH2�vC����\�J8H5 g«�p�PQn�եԸ��cN��IoU*�?Z�ݫ�����4ɵ�%�s�f�Ve��We����k=P�(�������^�0�o_�����4������zf���kS-ة���z��oz&�"g��-4�e���j/f�9��X���Z���S�y	Y���XW����-�ʞ�N�T�hRq�kC��A��M$1�����?�
MZx��L�+>�B���9!��U<�N30	Sp��-*dy�f+oe�2#-a���U'L����0�5��V\t�طT������)c)��+r��k&�"���a�Hk�`gN�j�PhH�˥�����צq�hd*0J�
�bp\�u�[�cvO�|�BBj���uc���G�� ƅۉ9(�WgA#�թ��N�ݳӪ?�-GcYĩљX�6��@Y�<�abUd��s�d\�UA�01����|�A	�d�Y�	�N@��I@E�9���>��X���J�ā���H&�A�QdQ6�=M����qJlRL�"R�/�,��/e*b�ż5y	�% 4E�qe,҅KU�3�,۶��Ҥ�����S�	U����h*u'oL��D=�`�E�S���Z@J/�oKiz�}�Q��3��A�Z:<p�ǫ\������]�x0�*u�H����K<N������G�K�L���պ%?�u����c�#��g>i��P��G�����<��f�H$�C��r���^���1"��Su_�Ӏc�A�Áx�vz� ��ܖ�M�h1�³l����/�::<ѵ��AHdg�n��!�	�(��sߕ1�4���{b�G�>�S���vM�"4�O��d}����qjvS5�RAe�	s_�=EI�\�j���~�Y��W�� ��ר��%A�|�daG ��|P�@���ap������ �]<�κ����y��_��@�� 1H�BB�`����<������ E����n7�h4�{鉶�Hq"4���?��n��+f�����8�\���W�d�B�MC��*m�0Y��&�
~ .Gh����@���X2�"��i�S�t5l��F,��3_ͼ�X;�ʮ+ǋ��L����}���Y���]�Ϯ���P�OJoe�rN�h�XZ�-A���O-C9�6�����Q�q�s�y��2�XAh�ۡ��z�֠k	'&Q��� ��'R3m���Zdd�ơdG�RBC���_�Z�%dg;x�H1Z�mo��]ES��gCx���%/C|ԺOJn �͘���$r=|�����;�Öj��������bf[�Ң���Ҟ��Bq�U2�����kf.����!���V�ھ*�C<�؇ �Lr!b~��w�f��f9P����W����׮�'.k��<az�����}@���'��&��m.� az����s���֖��d��(��, )����م! 'i�f��L1�x�pD��iv�T;�vy��]l	٧`-x�$��3�؍���~����Fa�B���҃����פ;�S��z�;+Ε�u�J�r[>:r��<]�Ǘ���cՅ��|�i�JQ4St��oe�`e����A�&˞G'�!��3\C��!o�{�N���lwkI�ip�����$$8�F�RA�xl&q�/Aa�˸���7{�Cp�q��q��BS$���.��&b�yv0���5�_���]
�Wq	�s �]�LܼP�Ci�"*��>�v�!e��r��P�L�ަ�@DZ����K���[�ӳ%4��2�E��;K�/�#^E"��'��b��': ���<����L�[Pq��~|�&1ZU�2f�t��W� J+|�Uſ&Ͱ�(��/PD�o�x�q
�=r;���K�-���%�/!�w��M۰:���-W:^�5����ߨ����[�'��Ay።�l��iԮ���������­�o��1�s�'`^S���uZ*Ba��P���Ŏ�L%T�jijH���0��+�{��!Y���N]i����Q@ϋp�����hrB �������LTef6�Љ2{ؼ���Q�����c�$T�b���¨�pc"�;Ԅb� TeX�ٰ��xiA;�0��ia�D��:�6Mm��-�����U�_?o�� ay]�}x�v�N�<��[ ���4��F�zO.#T+�N^?�
�����!*�Ŗ.8�O�yK㾓�����_��=t�> 7	#�6r;2�SXЈ���'i��'�\�ç�ȁ�?X�Yzrt8nW��|D��6mC��@�J$\��;,C���Ռ���s�J�揕h�&a��2{��H��aW.�!�~q7N�]�d��S��w�;e�������L�]�/Q<0�vM���aCG�`w��w��ji7#�oG��4ؽS�%uy=��Q)ǼS[�K��t�����c8�[��U�0�AƑ��N��	-MF��R}�f�N�h���?m5�r[�E7��	X�&�[��c�q�Q��>�����3�_�������+yg�T)`�����fj�s`���[u+����9-]��	�fKzVYH<�L��Ԕe�|}V��QJ���mbKW�?!�W���4�-�����������G��3�91Z�j
]�iV�ɼ\)m�'(N)���FUG&Hg���dy�8�V��F$��3�QN��#��e͓����F��Β�O��CV�<�U�mZ�U�8�	�ӄ�}��2n�� \��נ��]����S�LXVx����L[�M�V

`��\0>p*=E����W�
�7���J�&����2�O�F�C<�l��L���_=O�f�oB@�"�f�1�<?�=�5/��
��
�}��GI)�Z���}!/��Q��.&Y/��#�**�B'����̸��Z]u��."��h�^����e�_��w�h���q� Bu@+��fy��~<�ۘ=�c�j�d=�C���&!h5�	L>֭�����ݧ	�*3���0X^�������X)&2����M���NG�i�<̮
Ĵy�^~FG\�����y�?�D�*��.{�[�!�<9�נK���Nګ��� Ͻ�]�I�2E����r����Y\���kR����6)$��.����J��- 'Qaϵl�8|�DW�~�����!gC#=�%0�p@i㛆²7�l��߳V)�`�B��9���8�M�Mx��3^�l�@ڜ�v ���:?3�wmU�����8�5Vןլ��[���7Ҵ��b�ˇ�����;%�A��g���h
d�6.��6uv�vS-Ai>�ƭ��Q����oR!�YFb�j�˖�RfaAL��Q@�J�.pY���iM-½�։sI����l������OO���K�#�#��ߴ~�]��8�yd����{�����_F͕@��tؼ�m��5�g����hWM���=�B���J�7dG]�&��ϴi�83�rv���b�(�l}�c���e�\��/b�;�ͯ�I�W�`"oٟ�y텋��f����r�bG�O��y����E��P��!�)q��׋���-|��W���{����[��1���UB�ܦ=s�]��^�@����ǍZ��3h�}^0�������O��r!w���*��=��;�@թ
%�^}ڽ$9x=��VCu�/�X5	j��m�I��ޖoP։2V���`n}�Mt�#s������ �XaI[�HYP����&�F�z�er�r}>�
�s98��x)2��Yl`zF��;�ޗκ����x��	~����j�� ��+?�#,c�F��p�̐�EDNR_��TkF�@����NWd���vߐ*�&�lp���}�:.����G��1�B���;v���J�a���M�>#b�!o� A��H�ɇ�3V�L6H�z/k�}q|�c���8��V.Z�}ew��?�9s�S���2�+=�W�	��=O�2�O&_K2?��<����z���p��$��s/��7U��N�;�S/Yߵ��(#q�mX��pJ�c/0���Y�}��M
ph�^�����F𒚽��N��F��/R�J~�ed	�E�c���t�Dd��,7�Fy��[iŻa�<i͂"��j��@-�}��3���bHQU־�l@�n%h��+�3���dK���H���&�:l��M��Z���_O�6"W�����Jv��7����4�#9R��tRI�pRW'b��v��m������).g�eu3����\hA!�m�|�O�����t�l��P�h3��+���H.	�;8Pj��)��y���\`ID��a�`�EȒ�d�M�h5����*?J/��[��� ��b���k�|�bM��2x�0S�D���I�6�[X�jٟ�d`/jY��E���1���Th���됊uUEó!��^ "e/�n��Nc��V���.��#�J�w���J�z��	��s_���5�HG��"��,�Qlwf�eC�#[�-L/�T�3(����C#��9 *U@���lj���[T�|x �Z2����
��u\JS
�/<��Y��Xܔ��������[}�! ���]���O5�v&9��^A���I['7!�� L�_�C����xVJuth)�&�Q�P��5JƱ�<C�M��*�RZk�`;���%B����t��B��� ��Q[[�af�Ŀ�WpH�N����qa��і�j����t�h�R2��߃��J��9B�0�{g��n��'�ق$������'���R�$���6:�!�p�8U�����,���0G�1��.��,�����g�XT��!V��7 4y�%��� Riw�R3 ���m���C��շ[���|��!��l�s&T{p_Nd����.��K@ɛ�� ���s���)�1׉⦊�o�Wa�����S�gƂ�t`hm �8_0__][�h��^{�^T�w�|N��Ƿ_�r�	T	n�1���r����D�'���C'�B4EF22�˻��_�9��{3!�e�1�$�]�k�u�o$浢�))ҖiE$a3]���~؄���d��0!�=�z~P<5���Rz%��ç��EsN��-�)~����[2K���}�v��*�6��ʝ��0�L������[�eL���#kC��:��������U�^d+��.�Rf�6�A`��K�*.��y(>��l�(�}ө�2A C$�Q���[�'+{��y��8:��?���?6I�?�5��kˉiV�dy�
�]�^��IÑ�`-��=�j��\��,Yp&�h�^�P��p�*���T1*�Q����^n�ma@$���l�8��=����ul=u��]qޑ�z�=J�V\i64�� @�'��JE����bmo{�
ܣ���@��F|~�K�]^��=j�|�[ �-{���f��9��H��aAe|�'�έ����{_`=j��gӀ*�����
Jb�!czJ��� xw/i�|�{7t2=F�Y���ꬨ}E�#�����o[ˆ��K���X�1<q���%��o�b��	 ��겫������!*�j^uQ�����>wp�>���J�bR@:
��v�b�xi���N����q҄�d�k?>B�����\��(�j��x����S�!\��\ N��/����z�d��/M����-�/�\�щ���Ð�|-䲗���:f8��q	��O��,�v��s�?��<�%���DXkּ�r9�������J�]��=����eb�<ϑ�����@W��m9;
-6o����A���S�q[ ���;���i^c��f�kӜ�p+YF(~��S��b>��7`�<[���z�6�h}�1�uŮ��| W�k/�C���N��y�v���o;�_��%��1��n.\)�p����}�ƖO�4�zQ�@�D*A.��㽰^9Dv@�º�1��8���pY�|C�<HS��֯<�� ���(R��Ӥ��)Ɔ��m�g��dV��p7Se�n���
�$H��>���q�!�][ V�C�5�M�Am��1��uQzp�X�Qݜ����T�eM�1���_?&�3�5����. �*h_զ���x�'�����᧸�s��4ߔ&��Gpq��ڢA�E�h;`[u�l� �v)��
x핚1��C�um�Q�����է�	��b# 	!�t藡��I�ѕ�F� =�1��r���_�Ȳ[�{�OlNd�} �zlȂ�ܞ?�a��c�'��d7
�# ��sQ�kk����4%t��S�[&����N�������{Ʈ�zJ���ǽ�E��7"�y�q�օ<:m�j�/�syԀkݪ�R��dJ)>������T��X^�	7f�,JF�IM�j%����^�-7+:��-�V��δJy�.�ў��j�fyxE�	G�^�a
����Xl�tLr���$N�Y�~i 1�Ϡ��vtH���fsŠ�%)�.�qި�9A�i�,�(C[Rn#�U�����Xa��#���㒂'��B*�s	�oH���k��7��ȥ�=���H6;�R����{���_���D��=-��x�*?;����%8���)Caؙ��F�	�xŕ#����񢷟��ޢJ
��]!�����F28�0{vL�;0*Ҁ�A�P�	�+��G
�B��1YV�J�Q���ꡎ��^1/W]§"���j�8�n���I���?�4m�G�f�K+@��7��	�4�e��[`�L��
� /8>��[�W醋:���?��d0{�u�)����i��ԯ��}���9'�U�;�!Y˒�me[r�aNj�K�⍍V���Tlj�lk��N�����xO��w�\�Aε�ɿ�^���|`��[Ҭ�ĸ$s���^Qt�_��ߥ���Rj:��M-��WMt֤�9�al���f>�~aX���|�g`iq�/.P�|�����m(���6<�����Zg\�)�_�%�^>V�
��ɲ'1x���"�\�PB'�'��NV��p��R���{�1(���oZz
�,EӒ���[jk�BW�~kj��H��q��&-�&��u�����k����MU:]?��2����s`�C�� >����:��X��?���4��a�\�q�$Զ�����Y��M9L�����X_ũ-"�9�*�U�p��s6,�a� �Y#��\���-d�y��Or�q�뚕3P�
������Q�	�u��8�͢]o:k�TR���)5-��B�ށ���`6p�S�fR�} �U@v}���1^j~��-:��ɤ��v}� �^��>�pe����ޑ6嘟U���~��\�رA��b�o��N.���wFM/`\�o�D�u�����{���s��D�e�,�Ez��F	�!�is��Z�7��w+���~	��c����H����HUڢ�aq��k\�
s�����ʈ���l&H�a%O�ğ�����3��!BAM^}�x�t�G�')֍*�)�N	����d{�#G���Q�-a�1�@��ο�Y-~�/���Y�S��kWR�`I�gc��8\<Ay*�@�s��Pp?JzD���2��wx�Wu�w ��?4����Nv�"; %x��>aĐ Mw���~v�0@�Rj�4��n����#����`�)2%� �4Hd"!���þ;��XI���J4�c.��3���&�8p����YJ�� ��)}ߵF��6���t@\�Dq��k̓�95f�M��c�Yk�0��=��㙂�=�^������o���(]�� օ��ꖩ�aT�ͬ��ۈ=љ���u`�N�*&c���B�[���yJ<�)��md{IJ�\���[i,��{ç�����Wѯ����$���6čQcS\{^܋;�+�&6Бy�&�+����s��#�2�J)ę��T�Fh	��������`. ��U��/��F�Wժ	���m�:WnD�v$�O/��aW׆��.յ(��m@�D�ȷ��":�����?�F�&�K��A%z_1TE	-���u\g��^a�}�5�o�W(o{�+im �Ew�6']�%��[��+��Ըm#%��碗Ո�(	���}�4P�+mw��C�����B��l����u֨5���y~>�"r�w%�� ��"��H48����r}��+��V�F{��I���m^��=��a�������&� -�����}H����쏘C���0�QO���o�^��|Y����TB�{+�WD�p7\��Fo4M��WĪ�sMXZ��;+9M��A.���I���	nΝ����|r�[6ᵧ۲�������yF7D�I���P�v�PVu�r����C����l|.;���O$�*��8Pvm!v�+D�u1�}qe�k,��m�-y�W:���Z^1�A�|��7��U
O��m�3���*߸��7�3��� A���?�w{ݝ�WNQ��皕XU��'\fr���ݴ ��	XN�^SC�%�}�eත���u̿<�W���+�6��� �Ec�!�y�v�J������"��t2W_d/��Ƿn:残�Lښ����nZ��$`1=M�\��4�����KS}�,�<��^�ћ�E��2b����`�sS����C��F��pG0��C�'���N��C����b�
1�zS�����#@zq� ]�%~C!$[��8�ʌ6|Q��J��6�� Qq����j���P���6�p$bn+��b����P+GNvQ}�m�R9V/���qp�	8�cT��U)(&�==���0��8f����F��nPm%-C���:s�� j{��T�	�Y�ܟ79��!>ӭ�ybT*��v&,���C�*L³�<��_U�-B���%c�XM$�8��*�l��1;�ͪ�cY��9O|}�p2��3��T�����qiN�,6�D�3'F����X�z.���e���i�R<�xM�C�9��;/?.G�_)Aw�3��c����޸�o"c��#N�s\v��'IMՖ:i�K���0daIV��MUҦD�E����^�)�¦�J�=�n��N���xoڵ�R����*���z�ո��j`��3eP{�h�� L�^B�/r�)(����kx)�m��
!"�`��qSf��7Ns(���w����(ƚ��9���Zn�(ցա��]�'�X�+^���_��"�����[��x|,y@!vi �|>�Tt��*q�=!wr�`�|,������O��8E�.s��=c�k�I0��g~�2���y�����"�u�y�T�6��{��3'W/�-�XB�R�=�Sx�!.R�̵f�A-d'�t#-e3|[�p���X*�(Ւ�2�D�#�_}*F�v_-3�r:�Vq#�����]�"�	ǈb�w��_\�!�r���K�U=���v����
���PclS��R�;\�٘IGo�M*�����Ǩd��(Ƣ@�K�����f����/��.\�.�{��H$���ƿ�&"�Z�K�#ʭ�e�k��ф<Y���H��R�I�}7;,�-:"��,�Z�Q� �
�ؕc�8�����>��q�DN2�YB	U��#-;LF�֞y������h�f�~;G-w���R����u�-"�gh13wd���>��U=�=�l������鋎Y#]_'�IKn,�gjp���A$%�Xy��{�4�q�s�Jo��e�y�s"8i�����?��K�����O�ׁ(��q�_T��]L��2Bey�����L�`��i/��Ì~��+�Qu6 |�3e} �8��8�L����RG��f��v:J��U?庄Uy&�v��7�,�=��I��r�zO!2�n�5��NH�}躒8)B4��E��繮��&�$t$�� {���W���ëc�,X	��i�p=Tl�6�#$KPk�Bd ���-�5�H��{��m��0���2>
������!8���dJ�S�i����dc����3E�{�8��@�l�o�s*��	�g);��m�3��/���ě(5b��%�j"gc#��O�spwsq%#�t�D�|+P%�6~dp�D�Q=Kv��k�V
i�Vgs���<V�}�i�����9����.g��C�El�/T<�(�":�V&��IMd���wr��X�4��R8S8������Y�2d��u��F@�x���Eղ�t����r�LEA�#�ͤ�Q����PZ9vQ����GLu-�C��v��앧������:h�%�]Įz3�A$Dd�)���x�d^	���R5�x��90��I��+�c�u�Y��_��ېv�j��U��S8k�I	}����H%�'8'qbh����x��sK8�U��UV�I�7#c��ۅ3��')O+��+��#��cc��F7����ȯe8m%r�L�/E����V�a�$��c�/7co��_��(�?9�,�֦��j#�"X�U1TƢ�5���֬
��h����{�aw�$�>�V�݁��@h���!Ua*�q�-��"3�J��5����c@|���8��@�{��-���v��c�m9�K��t��ϟ�_C辱�G�����G<��
WH���y?��j��_Q�$'���MwD:h�A�1d�Q ���!�2y�9�^A��Ql���aL�\�5�?��	���7x�fX�� L������K�l$�Gb�����"$��LhT�L(iИ �	6�N�ش�<� }�hgE-uH�y$�I��teU���F��&e��B�d�併�:�r��`,lce��my��k����.|^tf�Ug�Ġ�c���(���yZ���~w���'���� &Q��'��o��^�`ʂ���u��6�V�h[�������4�l��&s��u����F' f�@a�h/0:]WY�L������?1x���w�)�+W�q� !·���!ik�8�$D��7R�������[C1bAz��m�JzM	��yq��|�]u*�^{7�"�mA�X�qH�ޫZ� =��pv$�v:��X���Oh���*��� �֧�����A��4P1c]8��hD{Ø�̱���o�q�\�o�#p)0��4Q��;�ܦ̖*\�� o��4mZ��iG�梉Ds��)pH9T�+1e�իA����f������E��� S\�kO;���	���<5����.Rn�{�M����(.|�J��K�O����bM���R Ц=^��Y \�i ��D�>h���|��CՆ9�O��X+��D ��gA6���I R&B���X��D0���e����B�w�;e1�S?T�o��'6����Jۆ�=?͆#$��P�&�/a��gt�%��?�Y���&s���0����wͿ ��[5�L�^L�Y���\A���<1o*����p۶�hBj�!�zb��OPk��@�`9!g [3vsz��G���8���o���<�*���.bk80�"
P����7{ƴ�[�g��ۻ��a�H4�U�f�(��1;52�ɜm�9�I~5
̚�0���L����
N8��HÚ��ܝ�~��1�vZ�q>�V(i�\�� ��~�*�L'�w$�K?kxhϳnU�K�$�V��x���dB��Gٔ�)�a(���&��w��1$�PoKL&���DY썉 j���@f��X���>�^E��6o#g�T*p�1̮�
�Ic[��8Z]練h��{�8�y����T� /S't����;��_8��a����G��W$;��b�پ��^�OR��,&�������zW��. o�ܾ'�*3"ù����H���j���`�R�4h��9$#�������M��e�+�L�B�Mb�
�ZX��\{oP�����w�7��0��0Y2��AYQS_b��{`K�j�Q�J��Gq)�^fL�А?t��߄0������N����d��W�A�����KA8·��p2ח�1�'a�v��cW��A�(#0�8:;��� ״R�&>�R�;��Hx�d%�|�(R{瘼_���z����b���P����^8[�$�L� ��]:vH���Zu��k��;4=�ԙ������1�����Mo[[z�(F�h�z���4V�����GJK��� -n^���w^���l!f9;�7Yx���FA��m>��a�}��C�2�t�)���c��*0���Jс��KZl�_l~d���)1W��V���zq�1;R� �(CŴ�I�n	fB � S�v��|:z8mq�u�*,��߶�P�D����_)�ƣl#Z��������+��M7� �;C �T�"�#+�=�1<�[9ή�to���)"@}ē�d�s37L��~	Gڿy�nN����K��䶡au�/PѲß�0�m.�����XBV_@*ĺ&t
�W�3#��a�\�ONWh������D5��s�M�ʢC�w�}�H��ڗ�$-�ߘ9�7�ܿ�C�R��oiQ�f�.�H9ֶ-7��~���B_�L��D~���`��s)�}T\�a��_s�#�y�s�^/�$��A$��)#7�*ۙ8�����s~h�)^��+��ޠ�3�O���(%��1�w~�[�'�[�u!�4 ���*@��7�d"���N��	`�`�^��a�ᓇ6�4k�Ce�p$TY��v|��3b���av� ��j�r/$��A�������0Lw��a��\L!*7��de��5@��`_s!0.�mxO�B�(f�cϞ�N �����D�ɲ��O:�<}���5M�[uᦤUM˖G�g��3GΩ�S��'��{Eͬf��'v��e��2�/ќ�-S���q����O�L�l�[�_����.�,?R*��}4l���`j����E��>��HϩG�wŵk=5�=g�&E�I~� �;Yv4ՁrЪ
��V/wZs�q�j�N}�	d��mS��{r�g�\w�^���"�����9�E��;.�����ղ�1st.����]����4^�X��l��Ŭ�S�}ׄl,;(��$���/%��#�蓘�3��L���a+]�L�4��.����)y�?��p<	�*�$������~�:)�@XỌ�̮͋�d3�f.����#�
8����<�f:����#���6���݆�h��|l�ɿ�t~ש���
WV���f�^�Y�:C��`�,{�J*�
G�s�ZX��w�S�����~j]����
5[�	�F̨��i����T��82���§���^��V��-���v▇1/^�F�8�������\Ӫ�Nة0q�tL�+���ɘ�C�~mb2��X�g ���bl���M���;�|73�4�0D��A�N��,��Q5�G���4�LIUS�"�f!�kV�~_-zs��R_���0��MΞ�)hV�Fik��<��Q���%ɴ�P���BX?Y��A.3�mV���\���2[D��krA��6�����Bi��	�4͡���b&]�7�M��*p1�.rA'g��	Y$s�lw8A������y�Bθ	�Y�S#|��*G��Q$����U�x��'݁��Y���@��Z��-�'
�2ܸ����dS�n���ݐ܌|׉LB0��d���j���YU���� Ag��#�]l��T	�pmۦ���� 1_����K�n�L�c���FJ�w�'�_p������q )u�������n���я��+���vV��O&�Ζ�o�>�J�m8�4�`�DBדz�_�s$��"uF��¶-?k�b��Y�zX�?�E�8�_�Pp�2��n�ȕ�!��c��� ���q�2�f0��]�h��I���v1I_96�"�v%l�d ��]�
����7����d�k�aGc�85�3L� �.��+�J��:�Q�]�i�\���S�e EXĬ3����wN܃ܥ�S���{�v�r�I�k�|2��ds�f�	s~ߥ�.M N��"7���b�[t�u���W@\��K5N#�����|E��Vr�I4{up�%����?���i���0��z�O+Q��KRO���}�k�c\&_ab�"a@����m�ܓ���x�櫕�Z���b���R�I˷��3���nԘ�؍)��974���_��-����IX���V.���!o����Ώ����떂�����Bsd�=P��	��=�G�F��Ad�ܑ �Ǟ.�
���� �j�Nq�$���<	/��b��u�laup����e^e^��b�ӭ�K1��1W�au��0��$!���7�H��p��h�+�{����.�bh��q8�	f���a��*��P��U�@�"�h���a^�vDOJmp���Pފp�,]�@=��,�N�C�Q��]|�W\���ֆd|�
����R��&8�����?WdXuuL���8�a�����s+L���MЍ�n����֪�A�T�y/��[�-�刴�r�0=�Ď�Ȯv�~�Tܮ��:_B)�f�j�ݷ��9x�v�u�����qơ{�k�)l����ƀ�u��aP�
5�A�=���@9ہ��yX٢B�}��-���I9#����I�B�-r���]Jc��B��S*	�����j�/��E��9��D+�L{D�[���%�y�)�2R��RC��R��D�M�	T"�,���
�!|Y��s�75|�y5�t8t|7��<A�ޗ�f��7}� ;�~����A_+�g�K�(��H�E��M���g�C"��H(+��x>u���
c����Vh�
�~��%7��;U3��!e����O�AL~���YTbQq�,�ZA�y�Y�E����5�4_��'蚱�۹O��������cI$�o%[�# U=����z����\L�oaW��Ȍ�,� ;��94��m��9��V��x��5^���m�./��lC%ȹa['�4)Qc�d�T��w�E�ka\'����\�!\u3�s��<=<�r��t�0%���LR�߼zl ێ�L�o+��5F�W��W�S �SN#c���a�M����w�.��� ���&뮍��-R�� c����9�k�+t�!��CwRѡ�0O�ҥ�g�;�P��ш�7WX�[�M�mP�1���*�	<W��:W��;��^p���w����"�60����L�f!%�<T��R�p,VMt\����ǲ�AJ�S>!e�:5Ba�F"h���	���.�A�7Ka^��}�$��o��>9����|H$y[ț��6M:&[���Wj�FP0��B���J����@��Ory�Ū�.Km��#D�(�K9�G��\�N*�tǺ�bD? 0�զ�k �-_��r@�5�4��5���k��L<k���;e�`t���V��r.6qz'\EEm/V��h�s\�{Flޫp�*��ݺMM7�&����+`^�OW�ۋ)��v�_�7~w��Q$2�����eg�mͽc�r���uσDU��$.w3�a�����������p<�w�t�c?nO;Nг8���w��'���Q��YW`͉�%�T��P�p^�{b�C��� p��"��[���Mg∽�>x%3����fM����x�����L�[0D>�>��YɁ~���͑,&�/��ne��G�
�5�=���ϱC�J�Pxr�(��q��\DOy��m��u��>�{�ϖ�_�:7�� �c�p�����ýl�F�o��L�lp�yt�G�j�U��A����<��U��=𢼊zN1�!��Jo��Ѡ0+{rw)c\�n�m/ �Vv�.͝+���y�mW�/.:��#{XG
K�E9�z|��iˬ�>��˟�]�o@R�F��y��o�k�}?\P��00���G���B
��e��9�F���W�:����W��<s�_��\�R�.Qpn|�4H�_j-~��.F�V'�3�j�>��)G\ÖomH���簲q��4���{��7]��N�!����Z��!���R�Q?HST���"����ْ�)�cĥr��ɑ�c�4a����x�&�^Io�y� ��	��¯֐
s0[�r	�v�Ҁ)��*�Z�� L��j=�~��
I����(�Q�Zڼ���*�����rR-e/�X�$���nK"���y��Չ��H�@�b�G j'�h�s�4=������)��Os��h�t���T�<S-�}XU?%�i��;۩/�k�@��,,��Yj�Ǖj�*��h���6nh�~�H�w	�$h��L�? ���-�k|����:������zN-�h�R���IeS�u�X�֐�6;�զg/���]��mYSN2l�� �/"*�JxY)<�6����m��2?^=$���T�R=����l#�$�KV���u�K��L�� �㰁�/���\�h�!��hv�/�q�$�������<:����n��z�ո����z%Q��o�i�,�
��9��H��ܗ���[l|>��cO��l��uGA/|�]�v䉿�)���}]���y�S(�361����H�
~j0ϝ���F|>�]�B�Y�'8쥈6�43�|�q^�[{�?Vjg4�� ���Z�0��N
��Oy�ч�Z���ER}SO����J0!qڍ��c���� �;p猉w���Wt�g��Hjf�5��#(���S�-��u@cT����0r��5�(����m�B���7��iA'�;�FJ�{:�Xoj_w=��Xe��j��g�XӁ5��tk4��GrpX	���`�R�MO�o4Z1%0R�5Z��y��<�S6Xw��G\�K����"`�P�3��|���Ch�i_cBN�����`JJ �U���43��.g����X-�� �N�-�ƻ�?������s ��(
�EuG��b����h�pn��N�g��0�F�솚,g�~znld:�V�YA�Nuv���a�Ɔ�
(l���Gp5UmvCh�7����3�t�Re�5��@�����f�|�~��b�}Pp��a�ni�'ik���n�瑪�y�YF��˝���Y�5�̖�:�r,B�&���9�SWF+zvw�yc%鞱AMzn��/�*���u3G$n ֜� 2�S������,C�i���`;&Ee������׎�M����d�OV��A��]41^�H�?QpS0��*E7'�4����`�H]��@k���to��r�f�!��n���#���Z��ơY�LyG
�Sԑ��g�����bEIX�wBkn�6�한��m�[[��2Ź���H�#��i��ց-;�uP�!���&�f��^�9�:�*n��Z������+�@_�.N����r�E���/Z�@GI�tiD�(�.mZ�T?��A=y/3[Ǿ���'	8���K������_�]�ŬMyX&]U���2�Xw�R̱M
W.�O��W����ry��Ǉ��#�;�1�N�x�@0~�K���|{�Y�*3.�]������i��{ ̾MA��U�K���W�K�;`x��(���:�G0���6U�b2��YX��n�SG�@�(%��5s�|���kUZ��!	�� .%����V�K}��dI^��>4|#	kکa|bdc�P6��ڝuUe\վ1Yb�7d|W�bM�*h�̐9�}�9N�7i���d}^>S�U�B�Ab�]Ҷ�7+񼶑��&ַ}�.l���3��*He���^c���*!�6Sz#1��Ěa�'�@�?���S�'�a�z����Y��ن����!�m�$d� yM;%�g��_9e���'�X��lF@s�J: y����FC�,������ �����ir�Y���5��e�a�s�(�՞���~��f���X�6���qH��Æ�9��3��8�9:���b ��j����TP�`�l���l�6�[k�-�┷�OD&��I�²V�Γ�?��bca7}k��:�1~��J�sF�J\��m��R�-5��FEݪc�������'0�����~�ld!4�,Ͱ�i�Ю
�I�9�!z�5��]�O�x@0��M���y��q���%�ț�r�\{cӞWc��ޱ�-�S���.��"���PݷA@��,�F�T����^������jk��`��;#
D�h8�t3Ê�p��2��;�J�B7|�&�[�]�}���ǩ�9�{�����w�بV��p�'/��)�"���8y����c
?%���o�}�	���վ��J����7|��ɒC�Ŝ_���4�|��O�gl�����%��y@"A�?i60"�z��C�h�Z��K�oԔ{���@N���'��hAj�8�Z[(%!�{��?0�`1��
��b�o8��R��8+yG��N��e��VӼk(�jF?1�u� �hS�S*ci	\�yn�(��O�ll��>�.�k�ؽy1K>�?��S���o�@�^�,
џ���(���B\�4C�:W�O�i͚��+���#��%��3�Ѳh�RG:��4�K��N���=��y������{&�C�� . ���K �P����_�u��ms��A�]���x�%�y�� �t:����|?���+[2�K�y�Yd��th�h>*I%�D@'�ah��R�R���������ƥ�U����x�z���T`҆s�h&�B띍�i]e|��h2i�97:�:b.���{@��)����5_��	LFme|X�U���Uɂ�^S�d[��%7a����,D�5�!��`�g�Ȍ�F^�!s\ձ��Y0d9���9��q�g�'s}U��*����g���ѿ�Un��-"9
A,�����)�X��+֌t:A���nZ�����h	��4?f���a�fe=;Y,5S8�z$�Z��� ����ৰ ��BM=���<Bs����ر���MT�P�T���}�K�6!>e��h�3꺢��C�O'u]>�y�k����oɺ�b�iѢWL��7Iđ�a��+��V,Ť�&����%>��;�G���vaX�Al�p����8{_4��=�!�|�u��f��gg��L�WHɴ�nE{Qyy��;���\)P��N�uDE�<��iUKn��IZ����~�!G�袩sm^�0��Z]�����VWu��$g�Uc�L�rt��2�6c�Ф4�A�fy�#_������u�yVh�+���@���d)��� �}��ۼb��^�ϑ�>
�	��k8�,�.�Q�
�$�M�:<��B�v�ވ�.�m�������U�m��{����i���uݽ�RfM��*U4�����:�T#LO,a��'.m`P�c�#,P���+�ɕ��~(�ٖY�I
�����){k�#��'�R���I �Hk��O���'j{��'i}
�c�C�뻙̤qy�����ڤ7��/��
V�_��)o!��U$��{�1
��N�h��u�D���kR>�����_�$�;�d,�ۤP(;���M
�d��I��:%Q:�Q�����b����S����7.��'��1\�g�vy�?D+L���2?5�`���:g��s`t�Ԅ(�P��X���]@6T=b[�Cc��~�u{��ȖpfQ#�,�q�eM�� 7���)9�����L���a��(�NI2����!��36�� d)I�_�:e@�� �(�O)��pc��#�
`zv����/��2��"�b�@���.yu>Z�%�ZnX��`<l�g�=�3R�H�^����]X��z<�I����� 7��y������{�xjo-� p���r��'׎k�>5����K.B�5�ev�SFP��Q���hR�6���2^M�{�v��*�6?�+)�d�g�'*���,sF�g�"W�ִ=�j{���(C>��d$�(��ջ��
��:=(@�d,����/��@��4��i�eqȴ�y��EN����:��%��Ygk�񈺓5��ԧ����<,��	'���eN��c�k�4T^�lb�QG��́�-���A!��[u.Es��CZ��
I���4f�\�,Y��/��Ra�O�ϗ��8/���erxOU���t�(_��@A$l;�
`��!p5a�$gu�3:���n�ۮ�	FŤ� ���z 3B�2AT[���mѸb�,��v_�����nu���L�(���.�mLa)�a4{Ϡ�0ׯZDEa��a���2$�̎���Ѕ҈��h��F����+'N��*��V�gQ��\%P�� T(�#%Z�[��Cc��'��Ӯ�Y����l�ݯ�z-��"I��֠�.ƪ�F�	��P[9D�0��,������t������T�҂�ԒVD�3�t��κ�	�:&��},yp`���0NT��߱?H1��7=�+$R�5�S�|�2d�/g[�����ߵU���{��9�6�h�	\	��I2qAP���l�4�N�Gz:v�f!�n@o�NS8��~�[(Yx��M��m�-��q���̆k��R�'��ʫ�1��q� �R	EUF1�A����RJ���:��8�.�ի7yS
��b�BN�ւ���~R����Ɛݸ��n�`��L������H���q�"A�����J`+��Bx�ͩ���]�B<Dc�绸��,0�����d̰m8e�K[;������U82�C���^Ƃ��}�?��O�1Zl`�cZ�C�ڨ�0B;u"M�^N���m�z%IEiO��l7��E�k�mxxO�)G߉	��B�t��t�@�+x�}ћow�n�|�;�m���
��W���?n�P�N��fG��ޮ�����]/��6>��y���S^D	���^���L�q<a��/��k���?h��/����!���*E�
��������RY��y���S�\r��p�{�C)����-h���l)	�����k�	ǻ[�U���qtw�X�wn��z��5�fYW���i}0����ע�T���6�Mw��OIV}�ŝJY��:}�˾��g��C���UE��������a�,�:I�?�G���T��ҕ�e��u�)�WUЅ�Na&~�Zb�TU���Q������8�VD"����| d}~EUf�gX�@�c��C��X�gR�سWS�s5č�rq�*U�A���q�&*Z�\��u��Q����^(�Y%��V�ϫS�p��M�Z�Ö�w���W]��p
7��\�؛rZ��1{[BWQ{jH�y�׹Yj��D�!���F�N�O#�Q6N��V�#�h�"ʱ�}�������ڃ��BS}=��VN(:D?�?����L�0�+�:��l)=��&�_��ȝ	��v#��_E�MD�-.��ZS!���
�O�f#悬	��eU�2 sUɱ�h��2��d��K���t8Z��B��ר\T �؊����L7��ۃ1��&��|�]U߂���0S��GM�=we�h�.!�/����k����D�1�SKGh�f^��-�Y�ɿ�8j}ЅL��A���PkRLv-���,�������Ci�@�D�.X����r�	NISߠ�� ��� YIb�:�Q���=�`غ��&<����h��n�[�Q��4&aI��R�g�8���i�Z��n�~�z�w~Ђ�N��:�h7�I;Ǧh�A1~Y��h@�I�r<V�?0Q�g����%W�*��:�6=P���]<�:�9ޝw_�H ��I*9"��6Q�Y�"#���,$���ÜO?g��0���{�7�^T+�t��Ơ@��٧�v�!f1ࠟ���Y� jID��q��FSt�@�)�,�6g�Nx�Yx�����-���g�/�0����t-�2-T�O������z�V�_g��/�ؒK�v�aN{�����A,{�Y𸱦?x"��V�Y�Mɰ6�	���i��ݮ�������&����nk�����?�4�����>V����J�C:�?3l��@����^�	�����L�G���%Pq��Y�Q� �.�{�
�4F(��W��z�Gf�Z�DG4��m��#O�xEX���aK��v�����Dmoz,.��@9�p�B
�/=���7���(s�m��a�����"�I3� F��̋D�8<j�S)?�;����`�D���.���'Cr���� ��K�fSm�	�ՆY�N�_,�-���Rԛӭ�����n���ٳ]s&�"
縺{��nF☔������P�Z��Dd.K
��u��ԛ����Sn��ěr�Ri8 �-^��Ȼ�g�2�"��am��m$X�Eϐ�Ӑ�6�}��p}G��:qd�'lN�,뚀%K�j��kXo���[.�$�C�׿ �[���
����9��\���K�|r/�vK��I�l�����]P�T���	��'��x��*���ᨓw����݄<m����g��q:��&�����"���z:�Q��l_D�[�|'{�s�I� :z�e	v<X琩`���"kZm��<����� �d �4��K�*��+����**A�p
zZ�'s@�N�9Xg	|(*��~�+\�q��V+H��&j�دֹ�ϻ�E�{����h��wf!�p�өs�8�9(�;?���ug�B�O��Ǹc�&�t�'K:b!1�⢺!1�#�m��r��M�͂}����\�)H|�� ,��4\����ZUD����W�Q�j�GQ��1��@����!ak˫8a]�f*=�׉=�!�^�ئ��*!�&��d_�0DT�u��b\���j����̰ ���]>�c!�bȎ�U^xN�RKy�|��Pf����Ƨ��g��߆i�E9%z�E���?�(T�l�"�T�N���JK O��@��P�r@.��;����9{�� "5'�}9�Q���r�'m�^�J�d�Z<�ќv� �α�d<�����1���XZ�NWE:/��$VWnȭRFhL3{�w�)8���"���cAo@f�Ϥ�0|�=��zD6"V��vDv�B�fNƷ"P��b{Ium!�6�v`����K&0B��U�dZ3h����䗫�d���		8'�X��踙8zG���Vyp�d2b�_߇��W�[L��^�/|�����n=��F��E.�o��\�n�K=�/�=�Uj"���f�ǻ�t6�/k`���^9�XV���%4���M" �����`�!Wa�#t1E�G��o+T�	��N	ډ�5ՙ���'eCd���E�����}a��R9�كĠ������ �[�%�t�d,��`w���$[�j޺����[�U����[W���ɴ���9�?����j��]��te��LM�$��E�N>�籩X��n�e%ݻe+Nw�^O1�YPM˄�F���xQ��r�e'���Puq6d�}��OUŌ+3lȵ3� ��;��A�ۊb{��I�F�ҩm�:�A$+�A�)����A���ȩV��,D+���y�>���y�4�,�p���s�f���Y�|�o���\�@�y�����ȴ7�Pr�I(K�O�DA���c?�ַ�'pX����<�.m�W�����E�Q�e>Gx�~v��^CS6���u� ���!p��j��>�}A�j\)>��d��S�+�'T��
Yb}�v��E�"��S_�OL����NHLA��Mg��~�1��YzB0�6rN�)��m��n�^�?��ov�!�@(qd��<lpVD)i+��$�����6�PZ�,kS���zՖ��ˇ�q��݀ғi���+����Mue6&۽��J�|$WW��~�cw�bZĶ�S��,���6��W⨮Ϩ\���6'���}�XYw��uPG7b:����D\����l�u\�����C��$���}T_���g(�g8D	��=w�_(�y��t@?!�kvR�mn
G��rI���v��@��U�9�Y�����y)	�(�t� �䪛�Ɨ�ݕ� ..�H���}��������Ht�!������g����n�	�����`�P���������ת}�֋�4E�_j��$�\>W8Y$�g����v�o��&�S��(���<ai��ח��ʴ�,ѥ����I�iBU��m�p�u �� -��8�Oan8�|L�I_�9�j�ݺ�%�R��1x,�
�S&�Ό�ò���U��J�>;#���[�U��KS�r�R��	\X��-���[��f|C��QG���ýxO�ʑ����O����V�V坅�P<�5{+� wɀ(h!�R\������2|�w'A�H�q �&n��#z��+rā�����E���j���|���|�Av[�!�i!Z��V����-�ل�����#���t��\�<5��8a��5H�=�<�SO���<��`ŝ�yi��7�����6��i�H��?=�Ϥ����"{�ʫ��wPc��:��8��~�}�[вZ���)s�-�:�ĩ��?��u6��[`8�R������L�>uෳ�������%oŌףe� �+%����ؐ����	Jz9�XƧ�K���w��a)]��A(�U�ɋ@9��UO��B�Lpv�.?)�U�rR,Z7���)�V�ߴ�Q+R�`�lf�;p�i����*�j��?(�c3(T��0^jB��*��H��0V�]���d��0ـF�Q#���vDttZ��^
#= �x�r���0�̢��e8��gc\"���-un�k�u�z�8W���v e;~1�����ɻ��f��a����~�2�y��p�sèM�ڟF+����i-���ڷopVh���76�;�@��<�kΌ'���O��(%"B�l!׌��؇b� 1���w�����rr���rQ1V-C���|������7h덡 z����j�>��ZE%
p��)�����q���2�'8 |��k�x�Q�����%{��}. �y��&���o���n�XUh5�P٬�?@�h��IXxl�ނ�\��֫(�5M0u��O��Jd�����O��h�0�dk_d�k�I?����p���)��[>�q(���u�
I�gJ	M��ϯ����6�%ΰh4���/^�..��gl��E�ecdF/��y8!�ِ�#�O��>�|����
�<n�����<�r��r]���.���f��(p1-�؝��{�jZF�%Ua]�"9.��yN9�ɺ�����դ��-0��1Ge�!c���rKVV����%\��`SrnU��"@UG Z�X�4̓�p~5u��,��!�����s�SL�J#a��,��3�"�!M�lQ��r�os��vu~�ԏ*�F��s��i�3�	A�5G��kP[)�u@��z��3��&��Ko�@�F�#���TvZ΅ԝI;��ǲ�%ii�=�_M ڨ�y�Q�J�HpW���d�@�|ܹ���f�~/%JOr%.���0�s�C܊ɓ��h�L��VǪ��l��|����
����&B�"g/&_4Z$�w�St�C�B:XI�̐��l�Hg\^{Tq#v2�(
����H�E���-�/,����������|�1>0���]d�GS��;�^OP�҂ùCg�F1k:��F�9=�f*�_���v�Gj��y�`gM>�P��BjW()������W���QSo�,38�Y����^O|p4��p (��WJ�-����&%��8�v�ކ+�����y�!��]r����P��x�O"�1h�E���h�c���#��׬uƬ�iΏ4x�kf��G=�W7b���T�d��uQ�%/���RaL������хD";N����a����Oޭ�i�8��%���l�WH���(9��֞�L�@[��	��% 
�qj�#��lo��7�m���RE�� ��9�ys :	�=a&��7��G�v����|냑�R�E��6���-d�Kťԍ�̦�����v�o0Ž�V��]�����d��$�Þ���i��Wo>�㽬��Z�4�J�&��m���T�B߻[J���Ϛ#$�8ap*[�+�AM5k'i�"��N�3T�Z�����
��a_S��c
���R+��x]=§�/=��"I��ȳ$��ԂL]�)���N"���hp*��\�4����Km��;���	B>�֓V>�	K��ci� ���A0DN�=Љ��#
���M�Ͳ����1����ˀy�Yj��Cm{S�����#�p���'tz��Y��
?'ȅ'o�b�g�J�jƢYx��������/�d}���df�!������	7���N�h��7�|�t��h��ĪU����2M�ԛ5Qb�]�:��Z��ɿ\�(C�ʣ���	q(�"����Z��'7P@6Yj!��S���� ʒo43ψ�F6Q�i��������v^�,Ĺ��J�Ѵ+	���� POԯ0��!��������@�c3�m��p^%w�G;U�㜐ƹC��c�a��q�F�:�zS��O;@������9s��F�N_=���l�kA������CC�İ�h����ջ�bG
�b��cc����h<��m�2}i�=�.]_�vq�qE|qVi�c�q�߿��5�n��!n��`>˶�	pf�D�#��|%?���"f@�T�b&����3,7��ͣ�����]G�;o�w�� �� ���_W�f��F�.��Rgy*9�tK���3�ZV��8�7ūkH���W%rM��g�K�f�b�o<��cIs��1���A��� 1l��v=��D�,FdC~�mAx�$��c�0�U��z�����L��e7C:I
u�yd��G�;ϙ��@��h���L�H�H�O!�X�@�����`�K1VPt�q��U��<���W�w!/	��ejX��à���1��p �:,�Wa���ñ��-%����sW��:)c����a���O����k�cNM+#���/v4�}}&́���������il��9����x� .�:Yf�U�뀪����â��RVX
	��b	{r�^����(�(&�7��
Y%��Q�g������u	��d+r�}�~A��ŝ�\y�
V��\L�a���S��������;�jw�y���崒��^i�R{�O��4��A�%W�W{� �HK���x�z�| .-�Oy�=���q�׬3c�-����4�:�l����g�ۍ{��+g��8X�~+3���
�۫��+q`z�m�J�	�����4>��[�HW'Ư�
:ذޤ�� 4�+i��Pw�|���ZW�a�ъ-�W�=��d�z8_�w='@�9n!!"�_ M�	��Gٯ4vL�6�BWr�,�L���H��"����wQ1xe�O�}uJ �g���洜�d|V�������h�=�G�61�D�j�5�yB���\�6.����F��᥵���9�ҳ�;��T,\�1�=��A	��Ì��?��d��u�G��rk{�@�$��N랁���_"�6�	����5�%8-3�/*ZEЬ���f�7q{�5'�mL�\���i�y��+��U���=!9�[s���_��Zj�'H��Ò�Pz!tp�"P��	�?$��~PJ��		��G�$��5�$w�(}X�U�gՅ���.����X<+��ی;p�	��ݍ�j �ajd/�����8� ����˿V�{\5� ᥙo��fo'�>���ڔ<������C\�X0��h᱂�-�iw�-I�RT�o�x�v��	�-U
!����5o�R¢R��'�j8XٵͽO��a>殍_-�i���Q��\]w-���,��S
��T�*!���5
����!z]	�J�z޴���*�fNRCP���$�z:L���eAX�u����5��H�SH��_WVʘ4 �Hj5	�t�q9If�V��4Y8�!��D��q��� �P}�/�@��{Z w����y]��h��t�3�7etF�d��(��L�aG��Eu�hvZ�`i�N�߸�?�J��x��pQ[�=�p29���QOtR��8��2�u�
��v��	�_��t�8UA貓��U�[�P�S�`��{XTt/���S�Ҥ�i���H7K�c*qx�`)�&��vcR�_��'��*r�X-��CkV�5�GL�N��o�u�#W`����D��ZT��? iH2��eZмSTS�vP���.STp(Ș�'0[uʶ��j�e[��G��݁H������hl�b�s�\���۶GI� \9)ͧ��+����z��?��y���Y2O�dC_a�(������j)9{����=C�x����ә���t^�6rG��,�pKiC�њ�r�'�7�]h���8Д�Q�R��]�R2�v��~���,�`�D'B:���:=ǵ��V,�����5�v�������$�bF�'�I(��3e�� �G�{�75xm����1(��<`��|�Y/~g�8�%��6��?���!�禋�ؙX�����Ŵ4��"�+g�X)��C����R���4�ӂ�00�p���n�-������z��m�������ӛUVt(D�G�z�\�>��y��#:�����x;9�k��n˴��&�j>�"a�Psu��U��#��i���9ϣ�y������H��kV����K��2 �J]�e�ӳۖ�Bx-�QFE/cv��:�l�e��q�8Bu�C��
��X��[���g�����f�e,
"�|'��t�����I�[��u� *j�Ay��w\n-
��4����1�8�2֛���Ѩ~���L����4�!p�yaϠg������Q$SA��#��a	.r`3��6!L2��՚� �X*C��%O�x(y咓%Az�WWa��[Z_�l<��M��E��@ZT���[�$�@��U�H�uB��5�?y�p�����'׳�:M*��2m�up&g��٦�G��@���o�w�͋C�ɡ����Zݦ-p
{�������|�0��	���A�<����3�P��ւP��9U�:�݌h�/;D-ˈWϥp�:�g춐��q��Y.<�:���|��M�1|��	4���Y�g��%��������):�}4ף*�O�D����i�0+��i�ӈ!K����=�s��Lf�#Kɠ�'+��j�Cؑ�U;�އ��b*��%��S���º�}5`z�a��S;棾s��� ����uvg���߳�m�}l�y���O���b}bڑ����L��Ʊ�����\�����de�90���'�S@&<���h%&�섞&�Ak�/����~�b퟿h]�8X���H���]�]5���w{S#yw�$�,��l'x�X��hq��k:�Lj������/_O��p�h�lb�X�9<��b����[{�e��=�k��5hN�n^�Қ���@h���!���y�sWf�7����ʞ���)����sq�Dg#�J#B���"x^��ݻt�,�@���a�����:7�Z�wF�:�5�M՜�:J��{��(�Q��k6gN�q
[�u�u��DSw)��ϹJ8��l*��n"�e�U�f� h!�l7,O/�F��c���9�Q�hLt����پøF�2�ȶ���2�n�������/.�L}l��O�w�ƚ6�.}ǻ�F�Z�[�4�S%{^_LWa����C�/�
s�8M,��,��x�}����zN�����Mg��4_�z3�++wp��eIĵfP��(+�Ý�3T�=/��]�[���@���8��'���EX�Ĭ��A� |�&�V�zv"nD�V^��_�n��bX��d0�R ���j��ZMN�e��P��m�|k��U�0�b����dg%��+�cX;7�ܩuH5�?����#n�#|�|�y���:?�v]鷷�������h8����z�p����40�`�0��r�z��[�1బW?�%������45al��|9�t/~�zy�7k�oj��=J�(G=�d�JzbP��N�%:H��s��R�U�ie5�/�K4�k�'���xda�Z�)�$-���/�9-��\��u��f�v�FY�z}���z?� ��=�`@u:`;��,L(ߨ��?ψnT��ԋ�s�����$t��/֊�2���=���UG��ϭH��z�!0c�T !��}��8{H�94���� [�
~HG���L��{:	��`/�<E�՛��(6��ѥ�Vp�;��L����sD�ık�r.V^�GZ `�!l�RL'����Y���(�q ��Q5;�l<��P��HImp�N��]��9��y���^P�}��e��t�uIt �r�	��!���P�{_��[K)��;���xd�Y��
z[p���qb/���y�9��%q��5�q</���XDjo�4/���&C�`��"d`1.��~w�\�6�0R�Ͱ��$��ev.m�KP����~ı��+��F�]���*z�OA��7�BU�S�U�;�V���O�l��ϵ��+��$*{q}Z�5����1��&=��%��D�펔y��t��v��L�L��x���]i M�@�z�d�d�q��l�0y`��[,���}��+���pm��.'E�˪���<��߯C_�bV���G߭�ǔ>0_`�	}�=F}�[�w��,�99�pBi���i��<Z(���v<.�V��= ���}�R^�䦊\�\�����	������/_�gcb��
=�3����� ~}�-�Ђ�?��Ź�)af�*2�Ѡ�I��no��RA�+�-2Fr��n�11�T�wG�"�.=�*��#&W�+ь�v�*��o
O#���;����C��;LW��c�`ܟ����h?R~}|�e�,X�����4�$�����e���������M�]X��OPt #J�uE���?N��3�B2�}Lq�|Tk�"Xv�3V|(�{��ߖ9 ��ėn˱1�AR��1��	/\�����+�7�*g}��ewu��j�t!P��9������*�]8��
P��xw�M�I�"I�>ێ�� �=z?q�ٟ`嵉'��V�g���t��b�+�Y��i��ǻ	ň���;���[�~�	�BQ�L��:uV�s'+����H�CG�=��<Ϣ+ǁJ��ӊ��qu��t�C���y��~��(-Z��Qۧ�^l'>���9i�� �W����IC�z݇����\���4��[�J'�������m�����XD���54�Ndl`���hYʺ]T_�(��@�+}�)�p+V)�e��\b���z��7�� �w�{�,�p>����JI�do����� u$P����S����0�(���>�'9��cZh���
���S~(���wŢ���
���K�h�}��\�ov���HR�Ŵ���|�tcS�ɨ��gg8��g�l����������OQ����/�5��ܵ��w��T�K���p����R�_�5by�Z����Y�������iCK'S��Wd]d	�k$�����>���^͊"qy���F����f�5?�< �u��hI���9Y��J�w	M���*Vܒb���epJm��-�GлQIF�����k(S�� �4�x����6W��u+�>�~�	����ǫU���lz�Y��ތ�������	@��>UV�� bfC`���֗[�?Q�9����K���:�&�R`��}���[MC��l�ͦ0��:�o�t��/���JQ� d\���p�y��{V��V5T�dտ�=��pt�e��ms��6h��
�`�͊��3ͻ��$����,���@���?���H����6C���/������V��kq��I_:'�?�r6 <AMQ,�O ������T�x�M��o;����W�U?Ā���<�B�z� �c�>)n�	�/��,�G��w/���OOkS�č栦[5��l:?�7UH"x�_��V<+�`=�|��ޕ`�&I=�STj=nF�ëzhV�l�))5x&����?���e�0�K�M���uq��g�M�����7�~��R�7�'�!o�t�=N06�?��L����w����+��U�(��ɏୗ�jkwRv!AQ�ìq�ve'aσY��{�����I`�]!4��a��,����/�-q���r�ݲ;]��d���tFި!JQTG�]2
/��C��P��kx~����I?(2P��{��y	A��
`}a�1̛���
C2#6�5�E���t��yǇ-�n ��&I��+{�)�/}Ϳ�R���+O��dε�I:/kN��p�kd��$J����8�=ub���G��M�K�l!v����*�C�ۙ�
*OS9�7�_�#�*~��>���Nf�H��f_���Wvٺ�&�"+u�{cSS�.}z�4Sh#� Vl�T���S����^7m阸� �t�I�R��%BM��\h6���F�x���VY�ԛ�u��6(�Z]�C}�&����7}�_�K���+�c`3���D*������/�J�����V�F��#3���m���76)A�\�o�*�v)(	�+��#\O,�;~��Y�4	?Y�<�+t"���ё�n�7N���C�O#��Þ͉ь\�nW^�'�..�d�wY�n~��`/B�ug�@	�gn���:5�`��HX��2󶵥�]��N�^�oB��Ў0�	TR4\�r�Z�;8����Y�#V�_��h��Վ�F0�V0�Ȏܳ5��]36f�&����#54τ�q�(���ə��vZ�Pk���{����t}�ұ�|�MQ1�e�����ܩ@�6h��`+V�'�m+�3A���r�Ņ�r� uɠ> �ڐJ�k��,��rЧ��[<�S��R|^t�≖@	"LI�`AB�zT�k�kf���ٞ�kQ�e��>R,��9��J?�[{;-��3�,�w88�#�XR�ܻs����os�:x+���Q�u�.േ2�y�_�~����`d8d/Q)z`�u
r�P�����4��>p�0<x���6D�vs@׬J6�4E+�kQ�ڂ&_���֟���̩�jn�mHRP%�#g�g�,(�G�X	1��q3��[]��v�§T4�%�o�m�Ԍ�Y���?��J�뾘4A�kn���:�;.��}���Tr���F+�������cx����b���ྀxpd��섹[|HGb�����	�eb��&�:��%�k&)�N�_l� �*�9C������7��˼!�����&�+Ϡ�ʷW��Xi^��H�}��om��-��K�{�m�SP��Ρf�{��ϋd�o
��:j�����f����2��1A?\,/vm�/����T�'���rNI� k��H�8�hD��)���eby�\�-_��A��W]�:j#L����D�A��`3���P�V��'B��D�����"~0��NI���k�RFI�&y~�S�B�yK����)�V�˪�g�}����mC�2Zt��t�+�8oEr������f�0�Z���?�֞��;K��7n92�rֵW;(�^��KY�Zmw�H����?K���|�ka�*�v\��Va95\��Q- �f ��(¦[l38"�k��ɂ�&g�b�ǭ�2��:�xR�Q�F4Q��rJ�"�]���`���dc(�nǓ�u�\�6�Rc�o��`�~рhmK�~�R/���Qa�D<��q7c���~�zK.���k*'�N(Do��T���u	O�C��
�a`�!PS�t�ڏ�M68�2�l��N��$���Ύ�
	�yg.�70��i�!�8�Fc �U�c�"'��0�B�P'�Kh�c�l���S^�<��
Ye�������O����p=��Z�E���ƌ��IW�IdN��ߟGJ�Mi�b�4�In5d*��7���Ch?�7��p`|�8Kd\2�K9�0(<~/��2�iN�_	�����*�*��$eP�D vS����v�����z�,SPRU��	���^e�ۂ^s0�$X�ў(�r���&{ �A~�2��=>3������d�h�WZ����<o>�wa�ś��3©����lr��j��|�CJ��8����,�L���X�������vLD ��u� �`O�p���Qc�@Y󯟝��:L!K	0�ZG�w�����l������}ev!� ����e����z2�Ç���������q ҃'tP�� �ᤁе������kn����|���n�������m�)��]���"��ym��Kf�D��3���zR8�v�j�ph>������5L�����Е+�H&���l�8���{;F/�J�L�+Y�08ZN2�zA3<�C�A%?(aP�􇨷��}��U�<ey�r�铨}�Y��[��ʡ�J�R�H]�N�yʗ���4L�8�*�(.���� ���g��ѣ_]o�}��u-��;��*è��b���-S܂a�����%d�����	n��u�DT���
�k�VM��q)M�: ���筧��I���觩�!�"%]:-�I��S�O��/���|D2#6�~�:�\
c���m��er%�0�˵�a��>���p����%���Ʈ�
�%��Q�(Ӄ��<\���������p<�.x���S;�	݇��v x�M��{7K"d=�f<<��C�8H�>�G͎O[G����?^	 ���唌�������!�q�� @���
�6�=D�E���8m����
��Ҷ��'Bt�e�p��8E�n��H�t�H�.m)	x2N䴐�WαM�oε��Ҏ��(�����{c������U��� /����"�5;�j�_�����"�}�/��(��~��9җ-��VQ�c��q�������T�;�9[�a�w.���V�+�����f鞗vKA�e���Ҟ�߷�s�3���w�LCt�$�=�C]�,��ٲwI���B�Csiq�xF��/����FPj�D)rD�:YP����s��~u��t��V{y�6�E�P�>5f�),�(h �l���+�|�ar�k2��-���w�n�.���`�x�!w�s�����5��X'�ΰ6��1�;�Ϩ�w��O '���%�%2:�T�R!�[ebHTV%�^B	�VԘ1������9��9���M������SE�c�� ��r�B_���g$��Ԅ
��0K[�r��2�U@�ܒp!;�Gh��&i��(�1���r�H�S4��پ,��&K��Ӑ�g��Z�,{G��Fj��U8!Ct�8���(5�;��+��;��ɉ�C��7HʿC'u��T�]��w�c�����I-Y�l���a�g��ԧ>2�eޗ�p�|F�����k�;K�4*:LUc���yv ���GkP$R�����u<�	�1�>w���-F)˳��6��
�2�5�%���f�8{�R����9�Q�ƕc�]�rU��w#�I ��h��ɾ� Z*�s��Y��$�@U��cs˽��~�at�+Q���]$+��<�������.��Em��S�p�x�vu���f��a�C/}��h�40�f�F��J��1̓P��z�8��0+�´�-rfÕ����l�r]����\�J�U`�'ʪ�h���]��4t��9��(��������6Ȳ�&�&�	ٓ){P���.aY8y�s&G��"/��f�B��=�|�bt���VD�<;�#��;@��<�!',���L
Z��o@]�	k�Em���/��^��"� ��HH��1pE�F̹C�Re��y��b}U�Ѓ ��5�LuE!��C�a��G�����%���� �w�F���eؼlԔI�|\��1�٪�8�x�G��"?HmH���ÉwM9�%>���A�n��-NG��S�0�-�6�ꊮ<����1وh�m�A1�&yݽH��U')4X,m�2�H�
�C��R�L?����"���/�=B!�1z�?3%kkD��Q�q���G8wy�(�WP~��s�:`���Q����^�����!t�������G´k�$'�f_� ER�5H�ފ0a�t�<��l�A�a��N�}w�.	���U���p���L���>s��u(`��Q$w�bJ>C#v@׽Y2���tJ��{�"_r\U�]z��A�qH�L�ڃ���]�XF���Il�ӵ��q(v[k��}�rA�f08'BX�.�]M�K����U�CM(�.uJ"P�KR���a�'S���ߡR95"�D(k�Ǩ�6p�ҽEE(>
��܆�xEy��<��E���K��#�����RFz���?mQ��Zfl8�8��q�2��� ���U�$����������4j�I���#��^�ѼԸ���_*ۙ�}�ti��W�*&jab�>�/G�P�V�P S�LPD10?8 *.�e�Q��`���-R�⡵��O��*���Fxd_���R2��X�L�
˝v�,��g��
���Xb�P�Q����ɪh)����ӏBO��z����w�+���o�i�j�)�$(���05	��v�5-P,��e�R ����� ���x�Prcޖ��ݪSںo�� �38��į%��8iA���̑��і��
:r�mh���<D(8o��)m�=�:�gy����V��*�����}nE�l]w��� m�����ۮ�܏'�ֺ�U�5�:d���p�=U��rP�7w7$	&��x;�
۝�mf2ڧ�V���wg�x�8$x���
���	�F�{'�O��W��{�Dx /�T����7�~1-`^�Z��9�U�u"���3��V�8�o�l�iW�}�������?/��� ��ڂVǡ�Z8�\i�۴�'�|jĄp��g,�|�"��4T�>�ֻ Ǽ/6x�Zxv�h7�����K��-E���$�M�GmX�L���e��������i�?Q����_��Z���6��	#���a��̀�a����r�����7"L?��R+�|�a:�PRhE�)�r��~,ƌހ�(�Ӑ��:T��6gBXiJ�@0�J/����Q#?�����"I��=���3 �^	����U�����B�HVI(���T����D�9n'�P���R5�Qz��{l�+�X☿�!�i+ލ�Ǝ��gxl����͛�� ��LoKA���.�V�t�8-[���Wm���1���_AS�����Z�8s�)�����g	�|'/(��@��h!�:�p`����C��aE�����8Wg��[�_�N�x Fo�VC����$���I����&��P;zaG_��`m��E�}擉�er$�I�k;`ã��i�c���_乥C*P_���gKL-�+����P��շ����j*���8*@����������D6A�a�ɻWd����3p;���Ψe��Iv}����[5�V��ν�B��36�yB��.����U�^QO�+G��W6�q�^sAV�f��T�s_�M.o�4���(e�R��8���Z�|zW�k�#�)Z�S"R:6���ij�|qXP�L���\���tU���,�=����M &���� \�;�����~x��� �I8�.]�3y�����0-�	3���$>7�܉��UR���عǯj���d ����Cv���]���9)�
�E~����]�vD�������ޝnKWD�y r�;�#��\����g����M?9�%{b�)i I�
 e���h@ԡD�
j}�!���W�c���V��4�꾫��j�K�+�1P�V��� ���t/c�?1��r8�o�}d�yq�����h�qq�(�ϭ닿na�"n,7���+vkD<�t�����=��T�eИ�iyO��RM%��Q$W�C�Z��ڃ>�ȂՎNI�qI��TM�R�=��9��fκ��v
�i�XN�a�2zǌ#�t
���x܄���$��fG�h����E�g���x���d�u1C7�7Nh�ID �.�/�S�YDe��ծL�dP˲��|���5��Xޒ]���X����JC&��t��S��V�IB�ȺJ��Ԇ�c֮!��T�EJp�V�F#S�Ƴ�3�:4;�
/�M�k���HA]��1n�8�\�jŒV�G�{�!X�4n�t�S��/c�-�$?֭�ZAN��̬:�b��'X��+ �
=��SWš |���2!�o2��{m3�t�T޶N6n��B�{����,c�?�M>�\x9u߸�0��9KD����o�(qz�*M�޹���-���X&�������}��HA%k�v.��8EwX[�TX�'��ə_�Q5~��+˕���!����F��V�!�(�ҟ���ۨJ�ܞ�>��5�]�;:�~N�����o�(�i��n�@���n��H/��V��a���nlX���Q�V����2��t1񯧥��j��.8,����CsK��99$�$f�`���ٗ��Y�F(ȕ��6�f�z6���k�( �+?���Xv���k���zMs�s �:,|�kEpw׀��VR�G�(nf����tϢ	��b��aC:x�㠒���'�i_y0�1�l-���!TJ�ej=k����йL��i2
+�^�q_U�M۱����tn+���(�.d��1+�i:YV5�R1>zp���L���5(���ϗ�^<,����5_�;l���"���{"�a����r�jPJc��IiiԛX�����D��_y'� N���o{EP� 	=j�KuJ�?M��n2*�����Rp��1�5��'�)��bt��ǯ�e<aY="h�)2aJ��4Lto@�������1����(�����l�9LC`	��)O����A�t&%������#7�/+4`Ua�z�"&e����ܧ�,��� �Wy㷇1s~����_����ZqU'�=r�l�M����V�����{<L9������j���,j�0�ؚ?��u���~�'����K�8��@�u�k��c@��j�ۧ5E�^�4�P���st��#�Kg_"�}7Κ-|	S ���;`�\�G��Hڎ�4�B�n����/�U���q�d��հ������.��>4��G�zQ�n��$���a�i��Ϋ���~��{NI�u;�`�����O{U�g�{��7�LsFz��_8Xg.�d��_n;�I��&d�����QHȣ��
�,�� ��k�(ɒ��b��]q[���m�N)|.�EjC��u��'ks��)�"͆�<���!.��޼����q�e��e����KD�8;�
�U	��?3{ԍv��u}��e�~Y�I��Zn)�(�,	���o�������-���6V���ɔj&�	4�^�Bj�~������'�6oYt��g�7�#��Γ&�P:�y�Ab��f{5�r�:��,�R+h��8��;�5I�w��V�D-B��߻�����t)��!���W:���:g3��dm8�G>Vz��F ,z~�œ�����դ)���胞��s���A$��.R��r�0tW5�֋�N�d�&��q��!�:�Ŗy�o�:X��f���@e,YշH��7�o {oK�"�Y��L2��2���r���۞b���;��6	�����_*���a��%ȧgulh������9e��ѝsg���Mi�;҃�؂����o����0|2e�u���
4f9D�;D4 F1��9����R~&��4�ޝ�g���o �2���b�{sX����ϗ�S�4��]�k2M-��~�l����竝8G�T��kD�������#�&/�����Y��yȽ�tF�،�b� `�w�i�t;*n8ֻe����H1�!G��-97�I

В�轫�e��X��� �,\@�u���)X�����S��n���M��Y"i�.䑻����魣��� ��n��1��v��_̯��l�P{I�x��߈R�J�������=�����l�<��r�^nDw��=���� 9�)�R1����n�Bw��IQ(�����ty6�
:�_�k@��#���C��ӷe���r�7�S���~J�ɜ�ϝ�ű���V�zS������;���[#���X��:�b~����[� z|���Z�>��~�B6 Y.�~Ye���k:G�k���r�8��o��v�Ϊ����[$3ڌ\ě$X��ȼ'|IO����*ܫ�M�4F��1"x�y�d���|�É(iO]y|]L�l
��?HX�c�И[q���� �C�qTQ���~E�",�<ס,O�	��'P�z�'�Ӑ{]� �6(�9��V@K1:���o�O�$�m�燇�9�e*�����g��#�fTn/sf���B~wQF!��_��5 2��_�y�.��Z�N}e�zvi���p���p����α]�Ȏ����-�g ��;~���\�z�� ���z�7���m�I�������jT���$&��-<.��h�.�_��o�[�t�rN�6K�(">e�{Q0�*�iH2T�]t�D-��+���^�E�ԟ�X�Cp@�\!���>�t�N�����Z�n�Z�ߨ�E�4&���c�M&Ϸ�5?bm�D�th�y2�"zG�
�Z�fȨ�^o�IZ��y�%����L�-�z��0�%��AӖ�ޱcp�eg ���)�Z�j(�
�
˾�)Ht���q!��G���`���\��v��V��X7��|bꐀ�0��z�(l�io�?.c�Eʰ��F�o���E��)*7�k��]��<��9��-|��J-�ԋxӦ��IljZ>CD�;u�rzܡ~�ac+�����8D獵���S�􊔌`l8��^v��9���K�x:[j>l�j��7�>b۪E��@�M�c�x;�Y�p1�
uH_��i9�>���Z0jB��mC}��5q��a07Ȃ'�$���W�Λ���cgd��I�$�S���#�s�	��6j���)�t�"gV�z7e�a5x��҅��t�ه�	۔���l��O�O���V��öbΕ��\��f�Q\�yD�S�<365��e��/�|�QTG�KE�0���B�p�A��z����V�*=͑(]�hX�663u>Ԉ��2���H���:spI):�+8K��Vv���>q�ַ��[�(EƜ�����CT"��1~��\D���⳹�A৲����ll_����R��ڞ�3���	H�~Ռ���NH����M�FE.6Cx0y815��"�m).��j���{g�S�߅t�NlD9�Z��^cR�)}bb�=�rF�9)�Њy� �8`,/�'7����3�g4�����r
ް�F清kG�X�+B�Oս?�sw���
Z^�����h:\�c�_v�8q\�]N�)�r� "�.�Kf;O��q.ޚe�\��Ҿ��7�(Z"z�X��]�k������BXq�]*IE"(�-N�b=E��;�fD$���Y���K���A�Ƨ����(���O�����(׍t�w��ou��v���o�X�L"����m��tai�cy�x0��XN`�'°^����X���Τ��8ȴ�l�f�Te&
=��2���ļ���$tX,
j�%돝I��:��Ѡ����ޑ.J�1��(0#.�PR���b���?�������mg�V���	9�E3������G$�L$��lbJ�V�Ѝn�X~8o�yJ}/�.����!o IM�|E�£&��&)�94�f�jj��:����m��;��F􇺠���& /�y���:�js	.�He�n�f3c��#�U��� �0Oq��K����yZ&�F/��M�3Z��SuP�k�|P��<��an`]&X��
[�9��<%��g^�Ϣ�|�y9SKD&��v�������CR�UɶA�.������v�E1�}Kt��9<�'0�2�d��u�	�K;��s�-��2��ě/�M{�U�O&k�!ϊĖ)���]�8��|��Z�A�Dt5�{/o����d�)�ק�sG�f�>%X�8B�qg�e�ٻ?t��tI�p���F�	V��1��L�����Z+�H`�=	a��UD^i��q�"�����Ǻ�FS�)d���~X�M#�^?c((&��iN$�0�ڸ�J�.��� gY�a�8��ů~�����	f�CCW��du��%zA��F��<��͕Nwe_�#`��iQ�ш���?�i�$��շ���1�pM6�7���x$��*@-{�8���w����H�Q5��<:��h������Z]��\����Z�%��6J�M�!�M:�ם;k>�?z�z��?�Mn�K���%o>{�+��u��k�vRgw�<��� �L	�t��v]�K/�+��b�?�HX��T�{��ؽ��D;�癳h����QL�0ya��~cB��FbS9��+����O�8��̼Sz��Re�)G:��辿�@)�}O����&`l���J4Kd��Nlf&���t��^�剷(R쐬��^trЫ�<�VG��J�i+�q��c߬ķq�I	 ��8����������c~P
���T�l��|�]�*Y����e:����o�E�>����h����͠��΍Μ��J���w-ҎƋu ͮ��5��ҿS�h�SE��ԯq�3L `�R���M�;��ة�V��H�Rb6	-�3p��h�JXi ���iO'��;ǺL��WvO.���Ú*���*˔C���F���yGF5��?�}A��O̤Q�(��kB(A�aY��TY�QL���&@���"���m�_�~�ˀG�k�R�e15��C/��Jyw�9?8i44���@�St�@���R�a�m:����P�( vՖ^i�v������Y�sE��&�z���:�|�"�P���"�QEVo&B� %�\Q�g��y�����:'~��F���+�g�6���C7u���6�>�2p&�e�eta�OW7q�2�'�ۀ�QqU���A6�W�^��)��RP�&�f�^�w��p7-G�F�\�+����&
*��rE�+w�4 Ӽ*����C~W��R��=$Q��BiNܿWR�!��r�-?�<����O��~/�&9	�HڲY�FP�MxF"�>bL�Vմ;�z,�2=YL�X��J3�Í�N�-�jU��è$���}CIl�Ф�oċJ@�W[�j�7��=W�^Q��[��D\��n�8��1� @K@O�<uV�O���A����_��\�\�r?���ZQ�t��|["�d�7(�_S$z�b�XN?����GgD�K2l��+�v��+(d楕RT��b�6���DJ�W���Hwn2�/.*�B���*�X�,6}A�݀AɌ՚��Ő�~�J?D4dQ��z���s\Rs���E��k�P�g-&�m�%8��"-������$&n3������bJ]A��m.[D+�����`�`�W�F�������2��R��I��M�?TS�}���GT�����I���L���R4U͆o���;V$�$��:~��N����D_�U/��r������ֱ���1�4p�:y��p�����晼��3ڢƔ&�:���A��P�ꙑ.��jSYY�D�t$���m�^/�'W�d��$ؤ%�pWR壂\�gJ"�z��8����4�	���e@��)���-�$���,T�s��=��Nx�_^�P-�	.�#�h $�?�ѬĊ��%�Ԋ��0�P��#�s����t���.Vhfؕ1.�����Ȫ�k2(����z] ��}3�wLg H������,N�^��B�E��^��~AK�}�.SM�LU#8��X��Wċ^E#' ԍr���vΌ��|n���o�����T����C��b>u�ߚ{v�����G��v�C>���=N쩤m)mg-�Z�{�wt"�o���2b'.�''$:}?ܡ�g�e��ځ�<6�p�}�=�/����A�j@�xH�`
��u��mpҸ�*!�~;	V�'�(R�e�i�@p�hjh�!�R:Y	����]����3���N��>��M{*:���$�9N����� P
ֈY��pa���mdi~�/�JG~S]o`��>6�lC��{RR�E�:g::/�lLVУ��s8�q�7Ѣ��G�hբ= Ux�UlSG�u�)�����o�8e�?�����AX�o���삷����A?��Ȱ���M)m�{'*��ŖT�u������u�[QJ�0\vH�H%�,��i �"�a-/���UC��5�]>!��Tw�o��� l��
RxM�,�؋{��"��Qe�c�@� ��{ß#h v��H)�\�l!������n�7�1Za����KΡ����O�]d+]���e	��L�4��W��hp����Κ�\S�H.z@6[��^42j��Q}�b�Oac���<l��0�h�c�D�X���� i� �����٠��qd� �950)o=1@���l��UBϵx�\��-6�%=��5����Ρ�t�ʞ������Li﹩�@_�;g��SGy� ������>d0�uc4�A��\Y������қ4u�p�Sz�Z;�t�{��"�q��v�g<-.���T�޲s�]�g�c;I�lq���t!�w<:�|�=�r�Ҽ��;�B��̀uo^F�ў�N�Ј�]�!����k�  ��F�艌�p�Y��?j�e�/-�U��&��3��
|�#ޛcw���ً�J`il�5�����0SXnPŊ�}�fTρ��S�r�/ �L�<�� B�V/TR�̳}�L�V����
5�3�C�3�H�XI���3�+_z&2��.�
x}��7���T
�-�ˬ��f�['��Ӏ�\�J�.	�F_w�2��k�R]���An����ʁ�b�� �Ig,b�n ��DQ�5'�mm�K(nR���79E��Ǣ���
��`�q�9��`3H��`� E��ذ~s4}2���(>3��%U�ь�3�]��%�zL�3�ñ��济���H�n��)VIP$��F�G�I)�O���0�� ��z..eFtP~�LEDx��<Cb�=��_��^�wγ�t�2~�]����r<ݑ�cG�\%h�S�n�4���
�L[y��N4�]�5u!�&��&����j"}2�Y�I���m��%ó��1t�IJ.r��K�ªv��[�젥��E	V�G���Ȩ��t�����v���~�4����yQ��U�)��W��%�ot|�Y��+�L���p\���r9���.'�F����%Vs��33�����t{]�m>�\X:�B�n�neg��Ü��$~�4�[L�p��$����ᶧ�.��O����ښy�/4�V�΄S�` o��~�J�񐧂��;I��Iњ`U����5����c�s�9nz	�!�W*,��1ض�d�l��*��'�{ن�x�	N�kPM='����н$�X�wL��,�ɇ�w��Ϸ��P}Yҳ�}���m:6���"�,�M����VQi��f�g�A�٨�e%C2Rm��wnY��a?��B1�A�@~7E�ߝ��k[e	�u��m�Q�t��/H�����d"��Uo�A�{�R��|l��Y��EǊɶ��oG�@� Z:���h��Zp;��g|Ӊ]��y�����#`���U��Z�Ͼ�	pm�|�"5��꿺7.�{�E����p/��C�Ԟv(O��vn"鲡�7���l����g�&l�&3���Z�M��un��_���u�T�q�:��J�RL���7�����0ʈ;֊�l�X�;����k^���6��4���^}�T'lP�>X��V{����v\�g���R�ТM��G� ������|ܩq��XBC�$��v����ǟ�B���|s���O�D�wCb�(�&I�\v�"޺Q�@F�����L٦�j�}l�7�DDÊ���V�8J;���B1g��;nhQ��r���(���6h^�K`�0]�e����V?o�6�R�d7�ŵ1N �q�z����̣e�	��IV��{�Ӧ�Z"��L=�$��[*֎}���$��qJ�֛i����Ӕ����s���!����٧#�f�)����b�?v+R�m�*p~��[��;�I���8{'�W���,�����.nSbͯn�#!o����b$��Yrv�it��FF�O��[�_��G�Y�@�o����mn��4H��=p��1.`^��T��
3��g[� ևN�����	g�Ğf�1���[ꢷ����N�ꭓ�=��eם��7�k&�C�Ȑ-�����Q��o���(��~��V�� �׻j	�1��o�D���;~��ԀV�TA�߈5@��l�h�X���G/ͧ%F:q��c�y(��x�%,=�M���r���� �l\Q��:��
��P-���'ŻІ�[+�a.�����*���"�0�o��/�x�����Ư���(��}��C�Ŕ������+/�������]Xi��=�
�����K�н藭�������q���q=��8c�!l�����=���������$���K�I��C�L,n}���t��,�?�W�`'*r�0U�,�{� ��N��a�ާ�z�N�z�1��
9�>�������H�!9�ǀ{8�;�Ò�^��[۠�dÖ�]1�}Ou���tؠ$8��]�[���`_\����U6�@��0���F��5�ZF ��lG�#'A�"��S %�Yi�q�#� )���|��8��tl��4`�++Y���S�T���?P"a#4F[�ػ��~�C���oo�S;��62>Ӏ�R8:z)o�Z|��n�aY�]�*�6�`w��Y�qj}���5v�͞$m%��IYXQ��I��p��%ɀG���Q��%Վ�-�%�$]\�ʍW��/z��]��|�Z�^�o٠��O�u\�N����@�6�H�{�9���ڪ��ct��M���O/�䛥�^0O�����3�Q���_T_uF��c����o��J��ČUWy��[߿zRb��
ઽ��@�����޿B���v<��f�f)"��JU+�I?����3W����ɍ��SW;�،�����9C!*Q
s��ކ�����z˛��N��F� L�l|/o��O���-/5	���˭�Mb�(��'�9��[��}:��	'��5�#���W��e.��O�NF�MV����W=�	V\�f��y�Տ��/�ҕh[�f5 �m!��F���(�l6�8;ţ�����	��D����U�P�K$�-pAj^	��ʗ��i�Xaje�u�7I1�Ρ��K�
/��+b���X�k�Y'�|��{�w�m#9l �J�Mn�I.�1o��ߺ;ZF�wP��K1��v����������# �!��Ԗp�Y���АH��V�g%�<b"�4��PkW?A��c�x�	��>�1P�~lJ��ny{�JTˆW��g�I]S3;���o��g`��>�xZi�X�.J�@�lg̊���o�O ��	}Ҕ�t��&w]������lF<�Vv�R��v�yVc	Y�����TU��b4>��~���}f�U��I�rOс���<	Ťw�NR9H��":��t���@7���1�#��ľ�M����I���3�2���=�X����'����u9`�6���@pK��*Y�?�2v���PP�+�v�*��W�
���a=���v��:����1�Nd(���ڛ������5�ѩȃ����oJ�!�o�	$n�"(�]�6��J�b3]/��hH���M��gsX]���Xa�2xJ�1�]�׎���4�)��b�(N�_p�x\�IN�x{dB��B��֠}�n���;���q7.[]ҵ�u�L�G>Ӟ0y|B;{,R�>� ¹~�=]�TLH ����ఢ���l��a�$�pv�q�RU�G���ag���G�e�p�zj�$���j�`�a��=ϐt�T��tl��$���&� ���"Z&�����L����-���?ӯa�=�J�ws:wB�<�����\I�N $�?鵌X]{O�h-2k%�o�QH�PUܙdw.���;���4�a�m	�xԙ�־#�cj� ������������s�x~��b��(Uɡ-�!�|~��e���]�%�BA���R���dhĭG �D஌U�3���ꖋ�U6�@X�3AQa��x+�4D��S�K(.���|�˽"�w�����@D�J�$m�+��ާ�d�~���oUԎ�Bb��<�!���',�JF���|���@���]cu�b|��V����kV����������_�f�C��� ��1��3����(��B���P�[}(8����J-T�X����v^z7�j/����.�����b\赞�\s��-{�ԓp!�R����|PP�L�ܣ���ƝI+�;7��ECQ�c��Ӄ�F�0�������0�"fuI�@"��2�)I�pi%-\�/��˹�G�Zv�]� ����\�"�B&�k� ���*��3*i863-U^�H�i���lJ	?��gE{���l��"<�H	�+Ǌ�0�]�c/�ʾC���Y������Z�ڊ&@g�/����1���SW�e��7rUa[a-}�Ϋ�������3�9�%\X�޸1���ߴ��
Ç�a{�r\m�������;�t�TܓM�D���@X�mK_}"[%ϻ��D���1���{�!\�_��,�]78~cG�u��p)���L��].W5J��wu�"�<�am��	��u�[_*�|R�ND'��@�xlEy�@彚}:"��1�bup��x��^��#�y��\o��93䫇��6�� Sy(��o��(L�����q�u�:ˑsae�3wAI�B�����&�''nX�"zɗ!{-m�	[��9>�¡�X.ھ1��Ѐ<�F���>\��Ԏ��(�>�Ƥ�氩�tN:��jP�]��MA$DbĔ�G{FVA�:4���[Ȁ�&��U-�|��S���������|$j�4۩_�/��nڸ"��\|u���H�����4G���Zf��7�5�ڒFE0��T��YR]bR>D��H�OM�n���O�����]�+�r���x2e�F8CQz�ؤy 8ρ�c�e� N�ftT�^b���T���� H.�iM��1���I��h�Xm�v��ԲyMR��0z�zl�c�{�R�c^D̡��]�u����ƌ��x���Զ�'�e�9��gny��Y�۞�B��
�����F��8t0��+h;���TBΐ�'�nؾ��:�;����Y��e(�rK�3̌�M�5��M%����c?>M���F�T���I%�j�kY��>�dA��*Z�cG��B�ʈ:����LPn�����]uF��l�u?�Գi�2�/����	��5�x��пʜ7��m�]���"a�uY�R��2�z����P��en�_��8����3����G���d�'w�)�
��($�3�!E3�JY �mO��r������ԑ����G"��^DV:^��<��D޶���bA.t�@�(��t�φX)��A����W=�A(��K�����hWD�����g#�y�i0x���dYE��?��>�m��h	�(=\�
'�W~���Cb���4I�	�*�XQd���>�V�C��-����6�5���qf�<W`�@�Ne�>V�nG�R���ӕ�~������PMD��3�.�s����2�9����2djE=�:T�)MI�ߕ����Y&�p!4V#��Ya �eJ�Ɂ`�Eɋ��������$�V����|�q�Q̋�sD%�6wӦ�6�,�~?�,��Z~p/�Z� ���X�j�|�3!�9��˄��EJ��g����3k���>t�X˶�����]q��N�.������3���X~��,H{5!��7�H���
lL�p��S~�mR	SKrYZ}��>����o����5�c�Ѹ��B1.����V��pi���7U�I�C'윶-�JE���?�S�A�8�݋�4Բ�['ц�,��B�F���i��Ȁ�q*(��-���d*�@���}�8�����OH�&qI�b�/2W�;��3��rZ-��Q@���S�9{��Cs��3
^�3��ݾ4�s��PS�a�7,�9<��6YOr@�Cn��09j&Ö�[��즢�M��vVab�K��׫��z�[�Ǯ��W���)�X�}����D�k���O�0�xҟzD��p��n����3��n�y샫Tq�/��\!���}�� �ʵ��S���L��*=VW
�h��o��.C��{�=#a&}"��ٞw�bds�m[��޴���r�
n�� �Q����o�ue�Lj�;��|Ĭki�VN��w[c~����]Qa��<u���&�$��:�`������%	ѫ��'{=����`q֦w���	YW�`�{r>f�ܷ	�!QQ�0��|�wz&�������蔽Q�)�f��s�!���������l���5ÖM���0��S.�8�����	�8�|�fE�Շ����ˬ��*G����^l�c���j��O��![�;��g��V�]�?R��U���S$(��q���Р+p��!�*���<粿�Ԫ����a��zع�|߼��S�x�����>B�hz쮅qaIk��4�uSsX%0�]�G�;�\�ER1��Z�� "�*�'����u3� �՗�Y&�@]���Q�yM�pY�u ��(^�F��9��/��������n�@���_���)W�� ��u�<�쐴ez���1���Y.�6�r��u^%����BJ$���Ƹ  *��H�2��[:z��?|� �_<�ń���l��y7������3G2�e�E��K�i��̺�0O�ҹ0�����Ҁ�;�b�+N\�_����E5k��� �r秨�j�c5Q�z��(��`dGf�
4���w1!�m�(�[PlO�K3w�U-�����e%�W@����:��M^�5��h��>�͛;kW��S��8��p�d���f���X�}H��O��`�R�/���=�����$2~��JЮ��U%���'y��(e86��y��5�AU�f
�3�4����*.*����|�@������N��>u&�5�X�r7�ޛ��R�=�O\�؝��?7;�����j��A��� �ٚA�WIP����*���2�Щ�Z�:Į�i���MC1#��O~>rj�A4m�(�1��a�p��1�je�V��͋�X2Js^��P�o%����m�������V[������dfi,:v��f/{�ɢ�aacڧ���c�5�U�&(+E����'@!2�A-P@9:�!����g������1�?��&�]����s��ݐ�2�	��;B���2������;�(_������u�/X�Z𯎖���q{��d���C{]<�_#�0�-j�؉R�em���ꈾ��:m�*���"�l�#�����`�.���� A�p��S���b8��{ܜ�27�2�y��BI�o���=RG5������J��vOI�J7����B;�M}�ܞH���%&��ؒ͋\O��@J��7�dg_u>��ˁǴ/gN,�և�!�6�GI"i"gҤ+WX��
�'5��w�+�`P�Vפ9��،5ڶ;��,�^`?�>?�c���fr=��6�h�Ul�9��}��O��8E��q9إ���J�O�߆<.���O6�p�Ka�v�)�TdC���.L>ߖ�׻��Ԧ�3�y��$¤���aɔ �a:�pt�e�3D�+�U66N�{��``��
<��ӈ��O��t6�'���Ƈt-�<E|��u}��)AЍ�����d�~�0�5�,��)E��S�x=���|�!>�\��p���FQ{ig��HD@j���Kt2<�����N��)7��k�� �酠h��(]l_�Ofi�MjM�~.A=��^��zd��1�����H��j�sB�9�` �_'wR��{p�O�(�̊0��v���~垁+^��sK������k�Ƕ��@���E�9gK����m�� ���PX"_:,��!.��U�������59q
9���\b�K�W�$�jbW��	0[�1�È���ʱ�6z&�^�zH'xX=��dOI�u2*�:�ZO�u�.�ͣ��K^X�l��\tUCJ�7�=NS���
;;&�Z��W=����'�p��'ki�IU��,9�?�NH�/�
�'�|���V˵]�cߺf��Us�5T�	�eK6a�8�fX�-����sqt�
�/�ZJx
�y=+�ذr��oh���A�V�R�M;Í��T�>�G`�'�ETh0"(����cx��E���4b�a�@��B��>y���+r��ͺa���E\r�W�5D'Q�1?�ڴ�L��n�9�ui��֖�ʏR��-Ԉ�,�x!�����(�
p��M*���ذ<@ep����[���Rs��o��K�2[v'����f�d��ݷ��;�2 ����I���`r�:y�7�'��oW>UQ�M	���+r��*cݩ�/�|MI��|�`
�E{�g�^�U6��-�J���.��~ᩞ�T#�m�hLz1�q�D�|�}����c�,.w���1�����7C��yM'���9e��D�-
�Z�W�����~��"����CM�|I�#1�F5�Η6�h�