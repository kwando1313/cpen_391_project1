// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:18 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Dt5CNGS7XW8+T+Yl2mXy779EA4tIs2iW+EiZr2Z+ul2s8BuG8s1Zs9vckDsqmxwI
q4UD9nsDDdcjGBCtUJTFiFhQKAv4wWDEoR/H6k83wO+L25AHluP/Juh+pwLrkkmm
5psDafRGJf/cwoNS8ztD9PFZ38krmgfxBR7clYHmEYA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16048)
2XM3uo1u1JM57mHOXNN09/+ASINDEN5yCGYwOD8bBhhAj5NZd7E8ahFbyGhpdOev
ya5anYq55HNFp3jwGxpRGtUURBn8HdOSRD73sUo7PZY1AvHtZttp2bxN/eLPOlUk
o43i2+ImpsXJ08qrCKElqBAhG/Q7ASn3WLZEwWvK6CfxaYa1kfWB3XTUmuIuKFeQ
05XOMsDx5n14kDOQnbXlG4NtKPkGLeA2y//z9skZ8yQWXES4P+75AFBWCqeH/3P4
RvmIhS24bptoAqEZz0N67ss3gwzW278kfbcznRTZL1K+vor6muHBmlsK3HjikFWD
bwH+5KINVVMAOjc2IrtsBRPsooI65X5ar5ucHMV1rRijaFV4k7+lZGXKplBog7Qo
v6FyBTXowUW72AdNo6vdjijhobadcgmpQGOpDrdVrbgLmWVJTZsMviiqeQRuwTfn
3RLpMIarBGnDYFbfpK+C7md19v01XFgRUn5ZGh944JD6V/XU+64edrhQjNnbgckT
NZU1ETyqyxlDZufQNNFwth/Ophf7uxyH8AAtchHjW/wlbiZ+qrcw8kYujDhxPNQv
JY5g4dyRzXx/178bHgz/xtgQTCM8eL/7eUuDtamjGKcIX8Ef2RxcbZv10GWBcv+n
J2mYx1lxefaLy/PTGBGBjUTo1Wd/+MPUlt33q+6EFXdjBUOtaVulLLm3o4X6AnGp
pjrearu+kHoids6rE87DHFagX0F3uPXZXriicDRgtkfLeepPh17knYX+xMHB1NaM
M0WpoA9ag0c5YEAx3+Z/MMuEoaCe00oOaHAgoeOhZHnt/b7Si/uQnpscrZQFeahg
7zPG8L/+Y0Csupi7+qL/IUhpLeeJvJTGBZrskbiLcSEavddvEH8lE2oAUUPqKPRM
QiBTwEkCXAqX8UIvcvUNX4psk/8IdurAAPWVmdKguFDb4CNtML5afYQo3AYOdm+B
2qQnTG2QAHiJtT6RGxfWpNNKDFVsSWzat88A2G/k5sf3lbQgcifv3GhOAmuNx4fh
3jYXDGIZy39KFYl76UcLnzixGDawFStLVzK84jjOxein10QxojrISmgM8Z5U1OfT
BN4hLC1ZdrucSrXNl9WjHJRxN+3nZ2x/iOO8p7WOH2xn/NV6CJ5v8pUP0I3tjqDb
DevP2/rqEXT21bJ5zxH7jJ5Wc3GleltihwB+VKvrIjnpp6WtvnKENW2Jdjw1Hpgn
YX0J7QN1++aG5atBuLJsXJJBrFh5RGqZQnDg59UboBAaTFI7G2zaWlM/4MgjN+hQ
e2DrTf2k/H5K0Ux4XmqCMswcVBmDCxeT77nri3mpn5bfKx6bzuETzulzAkVHmY9L
xY7frRkpXGes2utMLtEWIawwij0Xq5+CZkavFuHw2kMho4asgVrvz98AolSrDK6k
/UsSsRozc4SuTnptuX0mbsPR0RazFgTNIjNWokryzjr/i3szoJ5Xf+S2lPVOCt9Y
yeQWCLr2Pw7348pXuuqQLJIQ4xcSFgsCTexl21wrEURA+1rTNOu/Wo7dQuAC2SZ0
mGzbnpGznp7l1rnsS5+NhLp3ZRo0UCZG3VprBlilIM0AQSlg+2TabuYCWUWd80WU
TwnqJMc4IQ82Z6rAh9JIbhVFJKI4znpvwsMPkmDzQ1ZCPW5rT7U7pwjhns7bS/7U
x2ZBlkDFfk37DrhsGmhEn57P73E8cyq87Phfx1yfXMyUmFKdHqtPvEGqJCj9jD4s
c5ADsNjdoVuSKidwvLYy1n+k1udArh4S3TO6I2Y5+ngjEy2Yg+qal6olBuzUZlnn
hEqMeHMpz/8mMycS3SJQRScq6+7TRxVCjuz5cgOThNFUJrfgdczFHdrZ2XPTwe8q
mgx4Fb3GEC1a4NWdwwgKxG6Oha4Yob8yNhxYqLEYdwbVZ3sCKyd9tvkLsSVEU8zU
/5lJdT1ur379ZdIr/2t4FWGYbo7fddLruoXgB94z2acZTMghEXY2DXuixVn1K8GT
SNJLr/SW5Lb8URjdRFcUvvZ0vYGv2H6zNu9cTQssyvFq2oNmgdIKFnJAUa23S3/y
am7r/43dt02AlCEaB0+qmE1qMfCheIZVorNxK9TueDhM6zaeX8u10GeVcMSt4wJ9
lYwoOUWNQQLMQBWDTm0nwjBALIphRrL+M2sjBM/xuEW6RPgPbLOQ9rCv4SMYg0g9
V9YqX3RJnom38hfNL8AkNESdIg0LOt1JX13k6uc5ZDMCHKMngtwo5PAJI239ksI/
L78qv4EPOFIwv2D4vZhEv4tydW+9iJlosJIqoSFsvxo9OHTqBTfxH/ZC47+mLEPk
YHF4txcDgw2a7eCYmB7sj+DIgkHgsBEfhbKJ8hKdUOavVlTHE9wIln52nNzYrFly
itG0CNKNI9GY32aEQRtSQe8H1PmGo0z08mNrciF30OUaacglrQuWNrz4n93uYPoL
Rn6xrt5A8nPxmNZL2NCtL70VoK3kavHPzrGsbQcuQ0VPiwikkliWOG2AYIAwJ2hu
8LS2qIFVD7Tez/4AYQKawcd2+Pvp5KGGQeAZlDv1FKJUxlrUF5qWt0nc3clAF4IW
+EvUIA/3rCN6o1AgT3Ah1317dgrQn6tHXeVzREIrfA7mIWG6hUlZpjV3/lmNc9uY
Ebdb8aG5fq15ZD0sPjxTpkLC5wf1g4xFxls4NMP9Lh/9wpVWKYAK0JP6rTghOztf
Jm2Ht4rnDM8KXLwVqztX87MII6u6qBsi7w6l2v+x/Pq6aHlI2LDcw3GK2GQqgQlv
8yYaZ5EzcnA94jl9ZX/bjAl8KgIPqbP4R9t9TpqmJvhTRMALnEu7EfaLLnXJKTWl
aORLoxFp0cb3XZcjJA2j2XG45M0OMdBKUvkllLOrgh+BFHJfWrxwIcYuf+JkQQiK
NdxZZIN+8YfJxgBeexPh8MRqETiWHcV8Inj4F5L6YhWLjJIJ+XctpsN2b6fv4AuV
hxuBzrpy1CrrH6rHWpMBKXvBUD1RmvH8+bmrwd1ZJxmhTHjl1LCUYkgc3EuYSTWJ
rCRxry3smzwl8uFqoa+Euk2RmgQdRfEVtzPEkiO/KYs+pXUEkrH/NISdR6GmcuFx
AJzPexAhIZyx/RGEY9xC5Wu3Z1gFOI8ubOtt1hvSoEzJn8VsRq9kxQInM7UaGoj2
wBjkCsfQwUOt5z2g3AsXovdKyt3Sx46mCRLR0qwqKXfpT9rqibiyjuZgD5CLROL2
fYQXVb+CW6b7MJJG+vb4I8yEKH07puXhuKYpFPXigyfMhG+o0Zfoh00KajAgxiG1
ncU9ME+CYrTtoCkYOpV6703VcJ4RdZM+tsjcwQ3eLsoY0UiWQvT1JZ1PKzMeg5+e
UAls6HaQDAV7DU6Al2eBlhSI+Lyx4C8OyaXLHfk9HsrhsjjBUzhV0LufVLJmCwik
7S1u22TrhLUje+pecWECLZTPM3QOu+SrsskLtqROAmWOEV+boNcQ2DfrMD5SzYXA
3nYVrY0121WVfzcrVyXZB1HuHIY3Wun3M9LvF+q89PRG6m8ZTwjPg6PiIfDrb2sn
PolbJIMYXZZlqwj//WAvCTFvTDWbqz2EU4/LxiymMUsCBy6cDY27g4MCQ/PNdjh5
lx/Bd4sOhYxVVs3/jHkOEG6cKqpgIzLn0UVgF0PucWmabHgPoKs6/TrNu2cwKjMD
MZQVwvrursm8YfZG7Gbqu+kUwv5CB83J7wjOZU+P2Z5L6f4pijjekrPAq+23iIjh
jVRTV4lWMdlMqTb+akN58VmwTIaVZIy6qL0bNpfPrJJqn8ZzVhOqkg+AyJ38F4nq
F7uSQvxUFWhwO/r0UKIT0AUYVvqtxV0RK7c+PiTPELMt+a7T89Yz8AIW6gB7DJQg
seK/GZ5Pb2w5YZWHud5Nmm/8I3ilHQtv4TS9Bz86acJFmOGHv06Y69/keOM627Gg
1MpnTQns3TujaLXKoUzGQemRBV32f3ImpYwVGoeHGt5+YuewpzfiSDDhb0OfItAw
L65m+L0xqxlshyrSofnImv3UMKjGm7dotGWOux6t328dwklnCJznIAYvNjD7BYFF
vi//dTx1eJ9oLMi1zJ+mlw6VK9Ozd37VC9Y24XDFn5ay8aQ9xM3GWLGUcQE9bfQk
MCoCCaaueCyXpwG9V+wztVNq8LJ/tG8Fg99APuC1kE4kpaimZKtn7utM6t+oTdOs
G1ERGPvhqd3mAPZbRpw6HV5yxnbkgVDPp0Ugmt81vWWYj4eRMnqhHs+mQFJa3f+v
JKw/M22fA/ipAZ56tyIYhc/PP+y+sM1iOw4K8XtXZMzBJjQwvRxj8gKc2aefrfnH
MM7hJ4IT4liwd/SYukYM3QOctIkwe7CQetPY4ywi5oKeXRhPmtAGam6mUBjMVe6T
5Q77Y1bWD/62Lc87pqpc+V/zfjCFxgCQLrSRCtNEiksM13s3o2vd4JY8q14bfpe6
e2D7W23FZYqfEG19r3DUDJLSxUiYEq86SdFADdO9Br+CH6oAIb29AZlbiNKk0dkk
AUlr+uAcqP2y4doG2hDwQsHWnLZJWsmwxYpTDEl8m8O12rZu8+r/xp6wViufpauD
1F21hg0A6Jzh1mawnZh71Rt8bqsOgy4dy5XUxFsXxzsQUdO+ugc4YturbJDCGEOC
OPYgjmtv0mq2+uiacXyfIzCeOub/w8TfhrVV4T7jXDNn+0dYexZjuuY8GFhYU1e/
HjkAcyVdHuVaMzTW+/PN1TctcCDnLhRvnyiNttJRwozo3cilaWvyzO9hskCwk2Z/
rA1lfGZ29eEjrAdF5t08wE9XmBoT+AqphDVhrP5YFrZYtLA/Zob3S5cdfkTtlS7P
idi3VjYr2YiSdSShjbTc51BxcJcqFxunmNpwNfaoLhsZ0oPeYvLBrqlmM9oRvkT+
uy5QnW/gaIcGX1iOBIrFQ6zO7laQLi6Xdp9YpdS2Uu16nwyRw0D60elHHgAJa9+I
MmPTGcl8vHkS85D1Fc3yfmerAfiFQSQTPNajBf+Sz8mb3GwqRNtySsUrTOBz1/a8
kEJPydRwArrWlKeJLTuhXhe3TMqpGEjm1j9Ph8EwubZXPVF2YUZoTGk/OCfNW49M
xN1JLazkq6TB1BtcelzRg60WseLbR67EkajQ7zmN9DkuBjgcKsdXIaAaZ9xDoFIo
ZhWok16diaNAJ/u2RDICWun0V9kUyanKgquSrqW3tHwihkwFA2XRcc0AitnrxWxl
Qxo+tBYoLWzBA+aYP2Y26WVULFlOY5GgZ7WxFwS8bmp1bEc6jR/UVFi13T21cDwP
mR7kcesSc76+NlM16sI2nK0+wXqvO9iOb0/cjOSRsILLGXSOf7NcwEuWjDGo/s5I
DXKjMegAEQtKjNZtvMGjyaqBREqwxr+NrVyKBTGxQoY7P1N7l0RFg7c956H37FgE
812DwMzObdNU3qMOXcJMGPcBWpl0oLKgKjWxeskSpuTKvTxJc2dIUbR+DZaMzYvE
3OxrwWGT+trBhlzmKL73RxI0ZY7XP/jh48kjrbtR0mLcG6ekLRrf3bKvGYnxk7kN
RtlACu6E/6jTv9E+t4WUK3atUTyZuCcjaUH4h7DLxh131iOUcRWfuJjkpwjM+2EO
ssTQN0vkwl5Kp6K4RVozyxgkCzeVfKgOB//A7khBM2cJR20+D6BYO+UNFRL2EISX
IBFYBSpMKj9K0Z8OznkHEzt36oOdrSIKck4CrUpLsZAjzS17rbwmVHptL8DDCXHD
2qAlfdN5xRX9m0xnXgTrtEsKBW7jg9Pgerl2O3VcZr6DHkCniHnzLE+f8AfGcRvl
FOhFlFs79Bo8j43SGE/k8Q/cIaVhnJFcHduWfEnujocPfO+h6ggVqI0G+xR+Q4GU
Zav23Ws07NUwInChYFYANlpciBRVxy5LpaquTmq+vIj9wWh+jNA4dsgKAkgC5GUZ
DwFpZcA2WUUcDQKcagQloEYWDFbXOGqnVGTsvao8NsRNaxqbuGbzo7t75hX+782+
KlB53cZVtVuqBqcopoQWFaLi5IE5WAgRhrnh3Ua4cx9GJMI9LFqavURu4RE3ZTgV
uuHOhInnQv5mu1Fd/5wWGFwIetp13INe+7CZi8HVhmracExS7w7fLT/L4wxrneP3
doUpopdGNBxpAMFR2ZnD+HiwzFLlMFkFXuWt2W2xP+Shvz2fPMJcRhtumUZ6woM8
BemVurMT8IvnEY6/Y4mHfbuAJLFDNu2zjwJTsD4eZMHPAP/igoIlvhMtYhlne9hk
1KnvR+s3G0uBsGqJihkgtXbL7mt0t/XjfVGuqWUzkNKNDXgPz7LKiGBJj6vsQLdC
EfAcLP4pO5RACKtXaHTFj9z8eLQaFyLIHQWx4TacCq6ZcvpigcdVWhugEjHtKvXO
DP2KWkyyIXVV6uVc3bj9RmnwL2xOV7RueP6lha7yDAMrECKF01BzJbG1ZRC4oCVl
ZD/MBo53hGamAyhlD06E7S1N7hH27bJ9VIK8zKhRKhrc3Lb1TY4hLs3YoUQLBH/a
BbWiyLbeF1Z7wpOcx11Ko9oeX+us+eyPg/HYTED6gryo2ClwWZhX3VIovlM91BQX
8O63U8dItCIpzkL/EuDM8UuEn8gAelRDgdp4OfqbT5T1O6bhRETqo7M+L3g3p9S3
zSwFApfhX7iCD5mfO8it5IRbpWR+uVBs+4JDx7wpUa6xoJVCoHYbXLIQ0UTPI4Nr
fpM97z5gjPf9kfZS9tdQ8CR3VPZ4+W2W3pbn6Fqha3m8Yy6B+ow/RII3f5utv4IK
qE2mPTHHDOC/1KBKCLVUIWO3xfRvhtAYxTHA3aL2YlfJxc+jC6F7HeMxEsiLeaAn
ylGyggry8eMyPPXzUpLGp0GcVYzrfipZpsUVZY/QDCb9RrJrvn/ZKwi4ZZV8O3ZI
kgc7wne4KtQ+Y9RPj2ELX16lLaxlgZ3lzTbZyZCBvcfqIAulkjYYsipiEIGeqLC0
oDzOoUW84shqHa108RFL26N4SQmEEWjTM4AvVH2yVtmgPg65hccz0CjIlzLJSAjv
qIOrruxEAaGloiRQYFI+Z8MmAjK8ly2HZjRAs4prr+VAoQnuM8yFKeOIGK3P9FZH
/t4VctcDECUAcinYSFEcK+Pc8Gf88PYrTJL/tsOrHsf8VH0W1tBQOQEV5mkB1jbY
+gGftK4JgLLntYxh+cYJ04vyvjcM1bZ9B9VKnokLnZFxCcLdenEgxSZeNF1/tfh1
q6DDwvRJI2zpcYty08z1UyCeo5CDpDg1UXjr6ZRAbCv5xbUo+8lVbdeqdlm/R9EK
zoREfJWn/DXiJEKfmoCp8o1/QKbi33XQPPcUArr0UIdwxMm1L0ZEBTWUhY7QXf5C
EPdxM9h7yDWhTd3pk8/Ouhh1UcRdPavW9l6dng7JdWjopXmwwKDcVsyxOHSyEHz8
wpJ5quDArvVW1J/uG46LtucyWG1VSmqKs8pNMakyy4OqtW7sI7KCkLdIioA/z3bY
Ahcp/CsabTZYchkpCxevRJU92TQ06HklmvOxLGvf4ggLteX6iCTLWQQRNrGd/PUD
Im6zfST47MuEgrSnTeE0RBvRHiO03wFYLn0TfyaDXqvlcZTe2kD7pAwMheKYHwnK
Fe6LD95YIjhqq7l/pgOvr4TGSsLziXz+nutbxfwHEhVzqYeu3MdxDPntJSNTGfmQ
qDJoinaSb1EqhenJWwdGs2WeYHn4L82wtzqXcN8SL+40cHODaYH+XdZ0unMxmCFi
WQzBGlqsAgwM+NQQzzSK2nZ2vms1xHf7Rc+oKaFnq4ejA9SsIq9i5bJIyoe9qYEJ
78nN5CozrB4ZACQ9Tk3nQIo7KS1hOgypDRttJxg5N2IPfQoHX2TVvu1qv8X7jKY0
JNOLGmBF99bTABNF1nFRq92E0LCwynYYDjN8CqVNMRbJf52+e+E8qvoszDRREqSl
C5QJBU3u1QQzwpqZ3cTtFQ7Fx32mlO27A5LCyAvOf10oNZGVgzLfkN5eDwdHLRxW
LCfZ0Z+8WozliEH6k45VCcSA07Efy9ly66qF6b9H35lC5rXtABKC4CKpvOmjjknB
wdqoZUctFOyMuow/Ij12qqutuPs7AQ/oXmN0kdEiBf7/81TspFBA7UiXmo/LeMlO
CJhrs1JVpHoOYxLSWGaIQMad1DHkrCmtMehNcNphXPahOYLSr/ZUPnQdyqPo1L1J
qw8gd/CRzK8esdNa4LM5r8fnrtmSSf/+k2AebuSpJN+mL8xf9Np00jDltUeUmfGK
wIgPS6TJRvzJhgZtOlmWhkkAOgMA1vVLF+rZHUg8w4d1N99DjhnXAOw5V23E7sTw
lmuQZYM/zfakd4JNqieTOlYbVfjuIyh0inOBMxwYgjqwE2K8zwrpT/r11OVdLYmZ
fn5dAmFkxBuVEClGwzlWzY0dMB+ojdrbM/q9M8E4P66E+D9U1ZLQyJ1HLdwTXoUU
E8M7j928W98KTBU7xj1a19e2gJYAO+yHTFW9dx0pU2yh7OImaA3t4CXQUbZVEnRp
zDhVkkknjefc6RdNGd2VkKTuBFUi96YF/+dd/R8zTfb//xMrrKhvHTv3HCYxKdPU
umDBSNIiG9bBlqbODsq/9TWYmSWABao1RFrxhiOgBcrD/cNZe0XPNmSRsXkhzJ1S
MRA8ezX0rZwf3owvG35pAbLF/W3iSnLdPsoayXC3QC/mOSPUiBk/JHwQPIuYgF1o
+/SnfH5SnYFXsAP2wwTF7xPolDjKcxl57eUKAdPp5lPnm77YExkH62lR8ZWJSspU
jUOqa6cWKfIhG2W0dZnw5217aWYV7EpMVPlcp2xZi9aQA3bcLOCpXKqvkoEp1Sfl
VHViqExdIzBFgkFwKXIjtC68RQeDJtCvEnc+fnBBI42BV01SHyciYR99Z8RanlwB
vVYkdCAecCI+OaQmkxbr12YV6UmH52eDEQZEhIo3Y2wjYkwS59vA/+Trj25D96S8
dN3YmWm/4EzwNBrpv4/YvnU1onr6/eia4zwSZayAYovsU7W48VOTV7tIR6bEYocj
QHlxRTW2Cn/zwj9gUvJy6ZgtroUzdko9P/vMIbL9TxRmOpLJ7ExsGvnUHoH7mdwf
Px21JCssHDBRWj7Q/YvI01GYI3MVHwnJo+mU3wdA0+xrxNZXfhvv+Yz+7qFICZVt
qRvfKwJpcDiGXTB25xOm8/6eblKjxwQASa8s17909Dw07ZnJr42nG1J63d3MeSMA
OW/F2rgM+z296Q2sw1tOctj1sxzDTlegrmSUnbjAY1EFSyK1AVCzGQIjptoUtQ57
TAQZS2tkMHbECScrlYLHkBWf8WLKTc4kIvuMa/tyFi+5j3lb1giF8s8FMugwq1DW
uIAMzAZC9sXLntCawoNgUMY0Zo6P/08qAe02CIvjnhWrKKnAz7kI847i09x8ffgt
NpXnlfDU2IzNSpC64E0JMRwwGEj+hHlo4nuM4Hm5mfPSBVFoO/apTu5CS86AGpUT
lW6YIY5D7KaHemGvIv+htM4kXLeTYZ0M/uRb5Rl8RiuzZHAXHSsT+2jfhHyuS0NX
lW/v6ej2LEjTD+Y/JgFPII/q42OvGNl5iARIswvIu70boEZuWeoBiUFfI4wRohH+
pW1WbTwyD9VBMZ7uJmTrpZ5QREEljKeTFFTgXSii2Lr1a97KB5vB6lrrlHIuEOdK
msJ+18rP8Am4wY+IMoy7zOHstRsXDm8EGTSMv8ArbfFicX2j0SxLu6XbWxC89g21
xka3UdlIPVcRe5W+l9E4tm1YSVqgpuvY+inj9LrY9R4UIYYg9ZNMvE3d1iB2e+g2
Ujpbm4qituEnr13LvJ8KoO2asRUADvB1RbAM0MMVnL/eDIcxUeqb0MxjScIsGZYm
T6h1m5deCpR+J6r5RMbe40V7gktQijRdtTdiZ4OJRWDClUx2T25phr+xSo+8IwJI
O9UVR5R/re9HKTEzk5w0VASQsNKGubmYMeYAxQ7RAKIQfePp9J5aPW+2hH3/YJSP
8MuWEuTCxvb7WFakQz76Hhln+K0TtNGGbiX3WTUeWLJPKeHz/xf7raX87irojKMw
Ssy3RtI2OWwD3flaotdLfHLQvJGCgufydXTv+48jLokdh9xmjnq49TtxSwwc1v+I
JtfM7hY4CoIcdlz8myvwel+cHC379bMVhSpIhZLspIN/rwFkRW9KJf6E5QgO8wzk
YgMVO5bIFtBgGy6AD8bkkVlH6Qx/q71YvtZH0zDvqqTU5Xe87B+Cixd1WBqi8QNL
gE4wey8KHUcOA+PoagNmOnyw4s8wdIbqi9wG3YR6wnLYLB2o5K2GMiIWb/6lDdix
DF0GFtYPcVK7/BK0ETiMkzT2QMByn/YGZUGu+oNsP0EQIkfnkjy9LrGUzTKdSrhb
LFCzfIUdRL135QTHNkyUGIsV1jr808Ak/DTrgWdE6QQecKsaJ8LBvZP0yAFxHr9f
YKeOsIWK7KlrBiNqfuj8olYEReLqVX/HSreg8wqdwgHMXCBpYph0Mhkvttv9508g
0yhqDxZ02SQqv9CLI9hb3w8ig5x8KCAPBjuWSwGFAg/ASc2QBdkW38HVNn/qYuKO
agWi1jYj47+j8xax2Lh/XrakRGBZnSIO/FvbFITf+lU/c7QnkMbMcyIxYQzJZs4C
r8WBluKBVsFQ1wRIZ2bqjDaZU1aOmN2Mb9syApCRCCVi4CxWvNKIk+2jsuTgDNXO
vZ68oqnu0jFCibfJNP4Km0mlxwqkXqlrY9I9yf2LzvSL/5jLvou67uDZh3+xoqHJ
Jr6orKhgVnP0twKRN88hPbgW929Bs5/kzzPLL+jxFJk97qHYHJ+or9T8jcTcRhXo
hWpzU1yw4kz3V8Q5aRifUMDlrsGuHmkBxj2cEMFLoq8mo3srgJCNRlKOxxno8bQa
aSWSH/DET8P4ECyCNw7kE7rXfOcusX/U/G54VOLdQ+eah/SHs6Nt5LfQjdsISx1w
m6nXSSkWSiG0GgquxMsFn4aTExfuSLgHTC5abcXHdm5KiIe/lncD+uj/4BkbN9xY
WLzwGpmA2hxjKGIEN/MSrOc58T5L47KQ1yeRaXk035787pGEZaUfC29vzSXhbYWU
c3F58tiOhvfXY8+5NVFMM+bepsH74JccFD/ZR68DpwjVqwxdVK4CEeIg+B8cF7g2
8YJ+gdFZf9ZZb7cbALcK/5mOgplO1GlcG7jo9N8HHCOu85wqWuo1Z8TgKU1K7Kq5
76Ir6IMBz/y06INJQRH8wUVoylrnluwD4oIrsIvRUza/qhVlmOdn09Z0zzohfNRm
vDuJK4wDmydZpqGZwdsYnph8Ua1/mZYCDrqF6b9mdtcSRZ9zSqpI/qCUM7c2j7J6
ujnT90vDwOmxbQ7mMCIU/91Z/BGACV0HwsAAFe/iITZ1LuqahTXDajync1IV5XM7
nUmwoyL5Yjwzz/EBf/mE3arxlFGn1nvpdc1r/rKyOy9nNFxoJ2p2s1JRDYKRRJNI
ohiQy2MuzZYzLCeCt7wiVBhmhYOeU8dMO64O+j/fnlJFKtL5/mGL8s5cSy/UBC1y
leEPX6SfWIY+GsItti3DSbu0OAwMsVQUTvZVDUgGOXx7RLmtmamgogq8jCPDbixT
gMA03v6g5OsUdqAQyI/1I80KH/F8idtqkjSVcvduuOYfDhtOTELpCARdnO3wvxH9
rx41x+GeJxdQDuuQYMfyc+mxvqiqquThe/do3I/sMsKQmxkxxA1bkYe4qykTBW4j
rKAx03t7asBlMVrzB1ZAz3gEXqFjqv5UHNZiZc5pEVdaGBJj2zkcXhjJ6u4l2YI9
Fuf0jToUarSMnx4AGcTCUM36gXldIbrWGjjI/I7OCNm1QcR6C33qHzGQ6SgHlIg4
z8xEPLFQxk6936Og5K4vdTG9oDZjOljKGlpHA7J556U6LvGGLCC5g2ToUM4Wv0jL
Z0YfIMqqs6fAdQ8Uve17ODW09vwYQMosLYf5dftaHLMsqzd9RyJd9a92ILZIXbGm
zc+7yfLH1Sgurm26Ig9jCNps+j1xVmjHjnMKY1HvSJY55EKLqbXK2cDMRFr+rGHJ
HRaHQTbTaRKIZxUKpSp2Zp+4pZ5hgExNgl1EnBGLUGdiS/XB5G6aIFcCmFlrJ/bx
XanbX04sv1qghPzgSajYv5FZgySKhdy7zO7nbv4lpbt/d05OtuI6opmALN2DA49r
EMhsF+l2BYWb2Zggt2e/p7hgveMnknlXOpZ7JaFRQNGdk0r4mgQrF7YaVAQBm8bY
bTIcvO+STSAyxtME+xgrPpI0NG4hYmKRQxd3oG7kcH2nz9fJqp0Wmjk6QqkhGfrz
b6agtsaOPsQaqdmtTTUVJ0Em3kX7RhLKMS5b6eAPHCZ6TK4qrUShRt+ZyYjFjseV
gKrjShq9j7c30QIXBIC52ZyHcQKpkUTq+Cixrd6ab/2/r8yT4blAzGPgYHyGkA6q
Ri/GuoumFbJCgncHPsDmZrBbMWPowBHbpRBsNQKlJ7uezxyjhEUBl8hx+3frpigs
uL4ElC94QKOdY4ZgdMTlhgRdc/AmJma5oH4Ohw7rzPjfYWeOZDRxNfCYtYrrNCzI
LrLcn64mVmSU/cXWU81iUBTrVQ3ECS+T7NwpBLcjBUyK8ZSB2MBIjKWLlHCP7eNK
S5VE3zLsY3lJkQcuzuSt3t1IBC9ZfksVnW793m8vRdJ/Vtzac84zPFFb9rICuvgM
HQWX+9u41zoF44hlEcn8TAgtpxBpsV6ykM6Zy0Lh2pXEc1v/QJtbkTarv/YUlQtD
FU9GxHmTzHf7snAjqPve3CUf9ER0ZrX2qLI3RQDywHZVjSQoNhs5B1+AGZON8f9X
uInpYDLoVpSIEvjlKk3QguAXGq2/0ZsPtB6bPo9Rybl95YSFQxdh7xQVwT+2bxGg
HvyBx2E8RFweufManU23gkGJXiJVQDkYhNvYqsoZddIDNgQd7PGl+01J1wQk85ni
WBOLyEQBTqqXif53tmkrc/QUzy8AqrRPdYDEXr49ZyQT9EYqX9yiqMJcCOue+Hcg
P4oUbVFuSdCJssgsMOzs8c+7hxE3ukE0qNZWnB/q8AtBtv536w0a6PPS4NYcQwqq
g8Ug3m3i/iPLk6y1xzC2HOdDIoQy/FYDExwz0cnEWlZcQiNxIszB/4lzBWg3Dopx
A+IAb6BR9vSOI1IkT+9+IGi9Bm8EnRyouHqfGfKssB44egWecPU4DUr9exI7n6lM
sYuAfq83/Adwp0QLshdlCxq6Np97QTyHwd9hMNT4o7mQmrZ8+IH5mcZFYow8glQG
JfpoK6JajewF1MNSJTjqeZ6XjkPa0XLGboHAGRYqyHaEN+2ficntIo80pLRpJBkO
gWWnOrc/Lbqd2i4L4p9s0Uo8KPbkqmHrVZKr/BeTQco41c/2swHK6qEhpQVOKn24
+3DJq3nNzDvDPnB5cvZnM2Wio5Uw1nmD2R5oVgcDahPF/cekYMictrYd5LGwpH1W
THQIwUOPNAy8+/Fl4ZGsc6HxfSGf0fN0sYjjjqea6QzXGLL4988Rgkxdlo6rztRC
BVXdycdkGBXztYmboyZFheprj3CZMzMK/3eokQJOs2+F8SeQQlIvXdVWOBEX7/za
blnWaDvnsOoYVtOipSVE4E2swZGNYIstbFFl/n/abpfZN7ZNy03y8bG0e+ePcsnb
S4/iMFHoQEor8hFGVrv+YCjt0Fjyvx+5nYEgApnG5kiddGYrcuGWXvFbPWAiUnRK
hKGDVYZi1CwV3uG/QxVXus8T+JcO6/XdZgvesz+FsBVElJ7dOg5KYTH+6s5hlZIZ
Qk/uqObjZ0+u1i/SwhiOD1sCC/0Dfnz/SEw2NmTwpav1qe1UsW4rz2ld7oV9qjCl
ju2M9JFRS5mDkgcHkEXjQnKhCi3JvdJ3IUGT6AtBWLNLECAC0WGUW9C5WyyU9/6w
64SDpwKePXulGAJOLztEQ6YUHgH87QjzPtFXCdAkqICQkHrZav9hvBTKA83TOppW
qfCq8Oaj7E5XIGQeGTl+bZblVml0DLdiRNThDPImeczhJSubaeVB3rF0YXBp3u8d
web8pd+JqZ1VdyQSxSDMoMDMueJGQmZRtxAlzko1Drl1adX6i7uwm1CYcCu3v/FZ
efa+j4K+RfZ8P9G8eg7lqnsaxdzo6/c92jFpLJsHlgPr9/a3G7xsW8GRNmcIrS92
dJqIRzhnmaV/06g7my5mPqyj1tQMR4hJr9GqgftS2yb55RGeO3rAQTaZSRPhqezl
6jtIuCjcxjjz98IZaZhP2w9BIkpsXYf0hm6vhAM8hs+HOqdvKREbNYPwNovo5W2Y
rhDOO9wAdBiozysKYxuez1+eWkC2YzfZgUogAEoWS0hMsww5tpa1JerCUggtUruy
6ag+SFA+b1iRDe4G1yWPIch9h8HvvBaxN875ZWVh1HQGZqnu3AQDpq/mgnEmuhcx
8pCMbtpEYTeB9jtwmep/1Uv+eE8mlK0DqZO0RgDkYOSrossgdWOmc6OygBEap/SS
u5dny0abFCeUSxvSGyDjRehiByEHA2vh1YWWav/rn7Fxdrvg2nFWKpRxNfL4mkid
zSdKQm7NCXi3avKlLgbvpz1Fpc6HN/XWA3YRBDnyha8LtXWOONG6zgo+Xt038Ylf
xyfTLlX1kSGeFKyxkhKxmk5vdCtVmSJ/UZ9b9Ol4wT1pfnokivI40gVhApULMnNy
8EMotyCvNFiuXYQpCIW24IK1LKXDogsPfTVImMj97D5YX/uL7mAiBbD3IFq3e7xb
KJJ1nBghEMaxS4NewpnrzF51RZ9d8o2eG02xHIg4YSa/xtJtzTOMtLbAwOSZ4nPh
A9+Ms55r+iEE3FxOIyFbmraXSharbeUxTvXVYQ9UfrcUcB+RxpYTm9nRpormQGAA
qK1VHuzOeo2WmoE+DP90/dwe3HeW7raOX83kt3Rd94u4hGPKkIbpbxTW0E70iWqR
F/vEUlCLacpYI59uS6KQ3UAWc2m976ATax+o6Ayu5o2WIPjr35U+DgvGqLDBt96k
WCLgeSsmrFc7RLOesjvt5GXzF04EWpaFucmxSYTokS8RI1V/INdFjQGA9DETXZo9
KtYRX28QVNlVihcvc+03iQAtgVjfsuHVaFqBfdbz+XfFqNcjDMkdsu6hF3U+XxDW
DtcnuIMx1A+9FXhWMLvxutYZugXFFZ8GlQL4pGTE5+P+c4Hrl1hcExplsn5tmsKN
cF+7oZWNFzfV2u0ifgDf4/nDZtlBQ4rfRRx+M5LkgRnXYsohrlwMcNdFx0fNK04W
OSx8C9Vc2TDXa24AhlNY43aTmQtTUR9tERbN73LKlUVc0oDCWpOl2YshfrQB8kmc
rnvMgjlGP17AcRIobNgF1BinjCat9uP+mJ8leTi4h2Z3IlJcHrAiR3RfwlJzhH9A
g5IDZN99copwGb89VWw3fQe851QXsSpborq9EDlVM9U4phb3a668XTQ8X0tlzKG6
N2GvAD7Zirl/y6+dQDnFHLTVq2lZVixAPsJUz6h9nf5WBMPsaMM19EqK5RWm05Uy
r9B00uDo9DxDxkrgCrpsg5rfZsLF5POpi0kdWuelPf5+M7WTbYqYPAhb6H5/kew6
U/H2kYuBwfb1rqrKJPbfDJ8savLnowEoPK3+Jtev4fvBMx+zBUsLAdu+l0kfNCGu
ldXCYLSBXw2QC/BNTyAr0/oqe4os6l4ZnoQ8GvqN9bQWnPAun6in44dQ+tQvEOKW
aUXHilkTEWcgbHdwV+W47cGnTgUfg1GgZa/iCQI+ZUOvqiI12Os3eswWlpp+43uo
MP8nsKLs2xpSVDW/WWepl+PwrBhOMKwQpJJnbYwcA8SVnByC8U3qeAJSmrGZlxLQ
Q+MMdpPsPnz/JhSYKxwLhSyCaSWsVlDzRmdMNnHE3juGr0TkYpSyNRoZW2aRTvpl
vYtUwDi7I7JtY4Sf/v4ovStNrN+c2flA4As70aGLJXxl3uxaOPf+IIT0GJ8VYl26
wAqT3JP+Wd9HAWO4+nFrWw5rTY//9/sS+AaWz1O/m8M4I1xsMv/NGoRHQrDTR30h
xPwq/gR5AOyUR8joxoQ8PWrOobhhfWKSqpykbjKO4qrIZSFPpbCbOv9KqfTsvSEG
GFB1o5hbIqayZKj5xHD40reSsqFnorWWLX0yrHYTZmOOAp2tHkoJ0j5hNXJR+fKf
/VCf9I3egiBlhV6mSng8qUw2oCySwRRz6eApYADh4rYZo5lHho1Xw1JKnO2quPpG
A3hbiZ1Vmc3n0n96GiTL37PJpG+cJMpsuK7ONinExwiY8/kLIBtDRANYLB5bVpLS
fmLWOP0s4W3knSk2bociTDsXetBxroGH9FarE0en9uYT2DybW73wcJsoi3J1KwGi
VLhmKiB6E36JOs0JgpeWIpqYg0O1xyfUy2fA/HxHfF9o+BWYfZV1fN0uuASKbD0F
3FYtqTMKCvhgn6aq5MSEfRAMWVEWnOsb7OCV1LiQ8jNw1tpomwBxFIGbhmqy3qjV
dC3tvuJk63SXjbtsokrcDucqcHejnrZvgWXobpK78Tft8qPexnGdnHLoJdH0Q26W
VrARDCX081OO1UeaTkP82eaEnn0+bTzvU4523bn6MXWCrxHoR7s/gnZcQOfsMYEQ
KbBg+DeurB3gTNvZ7AXwdudkv2vRkMTizf9ZV7e2ChlSDP8LvulFTKtgsbXH1XAB
hGNVP619JBdEm1lV0wy/6oXz9TWEZwYTMLd22+SjZFD8MQycdI2M2FSQl7GDmL0K
q4fuRW9aZ245qTiwHUQHS5EM30AMfZyzhvm1g3Qy7QSI762WMD/9siBjNjkiBMUO
ksPUffVTAByljVT8EixXRtifiqdtfWdUK7XWR1RmLMxkMm8AP+VYrG74fn4n76x/
OPOGUFTHbMlzAMl+yi+QWzUDL5V8V9WViprLFsX+EJJ52f+FesUe4un+CU02mTY+
2WotqWOFjREXGlJKNhmar1YD8exR6t/i5NMZhR1jgaN9vNhkxV5nkUkdSnga5xel
U9m8okox0h6eXdRYr1wIRWHj3P6SK+frdIL0njuFiX4gfr28vPVPnH2VN6skPUdf
toGyYsJXLwbbUSx1aFuk/tnzzaLndK8s4lMJiRWlUwyL2XpS6VplRYlRiRL4f8TK
Q3PpZV93gpPv00djy6c9C/V/AoNUa9e+zuyg95W4R1aDOJjL3DaL4RR5spLApese
5LtRT2HgRW+K8khTU5/N+IUvDlova21GrkzL1f/Am6d1RiiNl0xQ8pJoSom0RJN7
i5naqoXvmT/ZguDoXYYq7OQv2gi1ZJLI7oECCnRo6gEhnl/XiwrkdpkWHoeyGmFr
yO1M4jipwIHfiTzeS50ZUJ8yzG6eBlLGpRkjoMzLWCgLvt86DFz2X6BANVr/tyAd
lk2UvEJ0oQCYfOFfEcUVhBjMr/3UHZJ7q/+2Q5CdUTmG8Ys4G2Q53P0ZMtgoHkMI
PHBI+6jdExjCsTApLOa07xKMrAT0+HmqUjkEZQR9fUU/Ld/jLW21Npko3yIOUefx
D9OAjAmF273UN3lUh+jVsL4ZADuq/45lwEcsELX7GFU5PLJUn0NzCp5dybeuU012
Az5mQtKTaObzhdT7759hNgSQb3tcrVv71bax5t0j1NZrv5PLRD4adVwaevLGi6yC
d3DFBxrlzE0S+NkMMqNK/N9JuNxYMhL0Dxup7MLFPvIcpyddrOAEHffPH0QMNaUz
A0tPW8kVAbOn8n/eaptaDJPZb9LnUsOii94S0ixJSwBlfjJiy73BNuRRcV+JHoHg
jaGtI9k7nqZse4ruEFiX10aNfNlvgGttSyXsxJvHXgNdf28L+dssTxJLWTdeB1aC
PyWE1D1JSOw1IJApFgVp5Xl/sK5oRzAw0OkwieySN22JMrJQaD4te9lXzHDDpdAc
RorvDNdS1ASnytbczsirRzz7p+yza7qPwjZPwW87gjjM1TDDpul8XQ/r2gJikNcp
8ZO5AJRXEt31aGF8jH+d+hNfrdOvQqb1jhnYc3eQyOF0KFL7iOYohGkI/RTUOeB9
X0cOHrKpPdWeReQtVBU6DvM0i81KUXH7q3zHvZ7gK8xjdnroS2CuG+q3s5o94MW9
dwB/s5H6r53IQuJhFnui+nfufLpFAJgJke8Kb7oq3XX9M8OVizfR23/qIceXTY15
dbAvCRBL7hRKaW/cFh2ntY0BTFmckMComB9lzP5d4wZXnDLanDJ9TP9/1PpA+9AU
L8JJr5loxTFS4awnQxLNP2YfYKIHbYA11FlkvkfYO3gbiTdVEDB7REnHGsye+cF4
RYszgPp2OjD/VESiwrn0hglkETNIEFpQj3fXJFXNip4ZSk49XA14wiLLI0mGKE0u
R9lYAzOst4xCoHA4cJqEuImbx12iIC93eU957pCU3dmUrJKaB4NNiCi5wtdeui27
WlkSFQIiQa/0/3aIdoAV3YJx6yk09rfaeBZHJw/oZoCF4Fe0+stL23NIkh4I4zlK
3bEOFAul5wShBVp1J7AmCnrHI3/G4y36dqLBb2Ki3xrRkn1B4W2UMviBIM4qpdg9
ouV6Cxipin2txdTdLd79gm6hjc6GaN2ZTD9XFo7YM9aMnuLHp0GObt+PNMBUdIuN
vxTFnkyT8WG1sqjR2LDki9etrbuQpDSteLRaHcF+MhO2bmWz1IQW+vp10C1WWNWf
ARMoLhV5gMeohFl9UTFb+NmPDp7anJA1A+EtiP6vQ9Xfj75vF+moi4IVzkbdV2XY
ERuu4z9mVOfuPEuBE+l0ec2HADCFM8DmihrGyOWVJjM/tVWoR2/uzvsJK0Kevc7p
Y5oz/j6CXWg9wSGU5HcHt7RBxyZVXEfXTihJUY9PES/MmG4cH9WoaozhevLAEHNO
Sw73C2NxkgAtusEc60RW+VfNBedDe+djlYOLTQxaQIbi5Z9Kf75g1NgNHQkt3j5N
E1hnxTQ3Egze4PDsXXIiiygqMpXWmL+v3Yri3hBjApynO04eb5gyOkTEjQ0cz0II
GSL18FNSe0TFx0RzjCA2A1Equ2UuqyiW1GWBjyE457+bV/wphNQnNLnEwy+ChYfd
HJCoQXL3LMqfln3KY9iw9GiNCt7zKbTSiP0vpXsPkp1GX4Nh7Wv6ARsU2osFXCjO
Yxue83HvG7/66C3cejN+hm7mpqK0lfXQE4an/amknvPYxrDJFujk7VoVtxg7Uvgy
vwf4iRABnxniaWVd44Voh3+3Hrry4SFR+JIB9oqbH6GU8fcZc0Tpd71rVGXY/ZAb
xOKPrSHoiE3EGeLsfSKoXqCj5RsKr1H3ADCt9adFNSTnjSDT4FoWpgkgBzyOqtRG
HGMxW6HySZ+uL9M5NSCjFW1FJh2aK0hsQGOMzO+YNpKa8wm1/JwKzF7nSDz547Gh
ZR4UG7d8AnQzsr9epb+oeUR/SZJrnCKy94kYV9QA96hSfsstP+FTD0IUQwYdk3+a
tdNYxdaM9FIslXFzOsm9q7FxIiCHQfoqzVciqqvjUJBVEulf4qayLWMKHEW9bqKR
lWwsNIsRQxhMDBzUjuYlGE0WfHhxofwCWVt7r37yf08L3kXuyjwKEwATpgZcKA92
hZqW6JQWmWxLlH/4xnVzK2REEeh+XjHnFOSf70MAkU7pL+0IHmeO4uRDN5Q6NYYj
mjPzWopCdGqqzomf7nkm7mAqkY7McaphXsvf4mkXw7VWph9Y6yd4YLsqq8ufe9Er
fFX3qTqMskax79toJuMP6QJJL/w2n8WNhOJeVKHzqlzsGoQ6D8+qwR0EdpnUTY5P
Aod2CJriQ5faBgPi5V/zxRGotUI/BQKhSDCLBarJdxHQ5+sPHhs9eYdAR6NdNhMs
hJsnWI4vHlKDQ82LStqLuDOdGCyfCm07OrRvW5dAfRKQmFp/qFH3TgGcas80h6nI
vvPaYzuVHt1RXQBOCGAdksBDqKn8O1MVKkkotwa22gHAhcR4az+gOEYnGAtuyTt7
KWVulCUsuzukYRNCAXRXhpblX5d9RT54UGcjpOlzD+DDdjneFejAag39DlnZ2AIn
3SZTxFmozCtsYyetyi6wLZC9UF294oR/xORuPLHYOr2aOru3QIaybPSqzHdB3fI9
Dp8WV96Vlt/se+pJeNbnwsQlwCTJSBBScVXRY59lY2qtIJXSUfsthvp5AlHW62hY
wXcM8Tl5DsDbr3Xoo4StOzL/9281sxvb/6zXv3KRxwPneWkneXCTLd75IVgIKEuC
KrzwRmO6+cfl0e6BClDVckhKb5Y9PNzVK1PYBI+hk2EF/utWkDxN2Wq1mFy4NBCJ
fbVIrbYfTheOrP4CdX+75y92ZKptzmNbvd8Kg6dPrq9ZFnlbd0jvT4IzbPU4ixAH
g1mD2OAiFp86IwMZApKiVwDfn8/DTPPopix85GrPw842wWni6uZv3O+IjqktBV/z
9Yds18J4MRddKWyZR0IQV9b+OG054Nn7rUkdgbYz7PrhEsq9AC495WBnniLGodzd
u5C4dJ28n+FZKUspwg6iIhNwPMkWHwOWybXbySLgVeueaG4p+PlSKK0rsR36A6p1
2qvp9DoqG7S9lQ8rwmO6kuQqf33AMKKwZ4q9459h5kzFPiNHwXxMWZ/e4Tf/kIsw
up0z3WlP928N/WTTOVMWiGTKNsdmIbs3mUq5o5+eGbT6p6UucwdiBES522SEjEQd
f7wf8q5k1wsqn82db1AveakDO5NNg+w010vW+Dh/QrP1LiZvFIBnvnM8wqJ7yP9V
is6EFE5goUhDsdYucbD862PBDzVSAr73UQVOELmhmY+fpk1kkyecMwFvIJs5AaLi
4qBS0ih0XNquPtjj4gfuPKvpey48JqcsJf+sk3+mSVo9uv5KOXwtXgS9qbhgNC3x
jqHK460Lui3AKM8BdAhKvI92ofKbZnRKUk4AgFXd4fGlmsIrhHm0OS6sYmIS0HyG
jGKz4xbEqTcwvqHwaAKJIRufHX0CgMr0ehLPR6RCuTXlk+R5nYHawiX9zr2tBr5b
ViBxw0ZMSuxK4Mhis3bU3NTR3DI9Ujo0wAbFK47HgP6tPQQM3/2zGJBFRuG7exg2
Br4BYBkGV240/lXA1vKnU0vgSHwTssHkPWSl9ubtSIYR1y5jXi2y0G4pVtL+0B49
YKG+tArf0NuvsMKwwJMwVFrvwu/9pkpDXrnq1lQ7lyedefcHBG6dEwYPiCNss9kJ
7xAKmPAWVKqKj1jUggTAKBu1MAY4t78f2MC+x30mt4EdrTmB8mB5CBONJ7gAVdwY
BsceBu9Pwr/sJVUnA2n0WrPYL+sMl2KZoIngEMxjIJgh55mod8l1PPnA4aoK6c1T
l9X5L8uS71qGfIIMYQD7nJGC3CMV04rhyshPXtu+TcoJn2121KIkfqIGgIpTv+/H
RD+5v7oTUq1EJY4g+GcIqPksCwHJMFU03Im4ml2tHvU1SpBMM/ELgme9QgNhQSok
bRKc2Xa2cm/rIWuZU6vtHFCy5A+kJPF9/ejCQWBFnZyZDEoODEzcONRRV5C1/GzT
iFG9iz7HdnlSrHbFl49wbA==
`pragma protect end_protected
