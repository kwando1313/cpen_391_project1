// nios_system.v

// Generated using ACDS version 13.0sp1 232 at 2016.02.24.00:57:22

`timescale 1 ps / 1 ps
module nios_system (
		input  wire        clk_clk,                //             clk.clk
		input  wire        reset_reset_n,          //           reset.reset_n
		output wire [11:0] sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,          //                .ba
		output wire        sdram_wire_cas_n,       //                .cas_n
		output wire        sdram_wire_cke,         //                .cke
		output wire        sdram_wire_cs_n,        //                .cs_n
		inout  wire [15:0] sdram_wire_dq,          //                .dq
		output wire [1:0]  sdram_wire_dqm,         //                .dqm
		output wire        sdram_wire_ras_n,       //                .ras_n
		output wire        sdram_wire_we_n,        //                .we_n
		input  wire        io_acknowledge,         //              io.acknowledge
		input  wire        io_irq,                 //                .irq
		output wire [15:0] io_address,             //                .address
		output wire        io_bus_enable,          //                .bus_enable
		output wire [1:0]  io_byte_enable,         //                .byte_enable
		output wire        io_rw,                  //                .rw
		output wire [15:0] io_write_data,          //                .write_data
		input  wire [15:0] io_read_data,           //                .read_data
		input  wire        rs232_RXD,              //           rs232.RXD
		output wire        rs232_TXD,              //                .TXD
		input  wire [17:0] switches_export,        //        switches.export
		output wire [17:0] red_leds_export,        //        red_leds.export
		output wire [7:0]  green_leds_export,      //      green_leds.export
		inout  wire [7:0]  lcd_display_DATA,       //     lcd_display.DATA
		output wire        lcd_display_ON,         //                .ON
		output wire        lcd_display_BLON,       //                .BLON
		output wire        lcd_display_EN,         //                .EN
		output wire        lcd_display_RS,         //                .RS
		output wire        lcd_display_RW,         //                .RW
		output wire        sdram_clk_clk,          //       sdram_clk.clk
		input  wire [2:0]  push_buttons123_export, // push_buttons123.export
		output wire [7:0]  hex0_1_export,          //          hex0_1.export
		output wire [7:0]  hex2_3_export,          //          hex2_3.export
		output wire [7:0]  hex4_5_export,          //          hex4_5.export
		output wire [7:0]  hex6_7_export,          //          hex6_7.export
		inout  wire        sdcard_b_SD_cmd,        //          sdcard.b_SD_cmd
		inout  wire        sdcard_b_SD_dat,        //                .b_SD_dat
		inout  wire        sdcard_b_SD_dat3,       //                .b_SD_dat3
		output wire        sdcard_o_SD_clock       //                .o_SD_clock
	);

	wire          up_clocks_0_sys_clk_clk;                                                                                                       // up_clocks_0:sys_clk -> [Altera_UP_SD_Card_Avalon_Interface_0:i_clock, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:clk, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, addr_router:clk, addr_router_001:clk, addr_router_002:clk, amd_0:clk, amd_0_avalon_master_translator:clk, amd_0_avalon_master_translator_avalon_universal_master_0_agent:clk, amd_0_avalon_slave_0_translator:clk, amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:clk, amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, burst_adapter_003:clk, character_lcd_0:clk, character_lcd_0_avalon_lcd_slave_translator:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:clk, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_002:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_002:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_006:clk, cmd_xbar_mux_007:clk, cmd_xbar_mux_008:clk, cmd_xbar_mux_009:clk, cmd_xbar_mux_010:clk, cmd_xbar_mux_011:clk, cmd_xbar_mux_012:clk, cmd_xbar_mux_013:clk, cmd_xbar_mux_014:clk, cmd_xbar_mux_015:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, id_router_016:clk, id_router_017:clk, id_router_018:clk, irq_mapper:clk, jtag_uart_0:clk, jtag_uart_0_avalon_jtag_slave_translator:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter:clk, limiter_001:clk, new_sdram_controller_0:clk, new_sdram_controller_0_s1_translator:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, nios2_qsys_0:clk, nios2_qsys_0_data_master_translator:clk, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_instruction_master_translator:clk, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, onchip_memory2_0:clk, onchip_memory2_0_s1_translator:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:clk, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_0:clk, pio_0_s1_translator:clk, pio_0_s1_translator_avalon_universal_slave_0_agent:clk, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_1:clk, pio_1_s1_translator:clk, pio_1_s1_translator_avalon_universal_slave_0_agent:clk, pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_2:clk, pio_2_s1_translator:clk, pio_2_s1_translator_avalon_universal_slave_0_agent:clk, pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_3:clk, pio_3_s1_translator:clk, pio_3_s1_translator_avalon_universal_slave_0_agent:clk, pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_4:clk, pio_4_s1_translator:clk, pio_4_s1_translator_avalon_universal_slave_0_agent:clk, pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_5:clk, pio_5_s1_translator:clk, pio_5_s1_translator_avalon_universal_slave_0_agent:clk, pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_6:clk, pio_6_s1_translator:clk, pio_6_s1_translator_avalon_universal_slave_0_agent:clk, pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pio_7:clk, pio_7_s1_translator:clk, pio_7_s1_translator_avalon_universal_slave_0_agent:clk, pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rs232_0:clk, rs232_0_avalon_rs232_slave_translator:clk, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:clk, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_demux_016:clk, rsp_xbar_demux_017:clk, rsp_xbar_demux_018:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rsp_xbar_mux_002:clk, rst_controller:clk, rst_controller_002:clk, timer_0:clk, timer_0_s1_translator:clk, timer_0_s1_translator_avalon_universal_slave_0_agent:clk, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, timer_1:clk, timer_1_s1_translator:clk, timer_1_s1_translator_avalon_universal_slave_0_agent:clk, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, to_external_bus_bridge_0:clk, to_external_bus_bridge_0_avalon_slave_translator:clk, to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk, width_adapter_006:clk, width_adapter_007:clk, width_adapter_008:clk, width_adapter_009:clk, width_adapter_010:clk, width_adapter_011:clk, width_adapter_012:clk, width_adapter_013:clk, width_adapter_014:clk, width_adapter_015:clk]
	wire          nios2_qsys_0_instruction_master_waitrequest;                                                                                   // nios2_qsys_0_instruction_master_translator:av_waitrequest -> nios2_qsys_0:i_waitrequest
	wire   [26:0] nios2_qsys_0_instruction_master_address;                                                                                       // nios2_qsys_0:i_address -> nios2_qsys_0_instruction_master_translator:av_address
	wire          nios2_qsys_0_instruction_master_read;                                                                                          // nios2_qsys_0:i_read -> nios2_qsys_0_instruction_master_translator:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_readdata;                                                                                      // nios2_qsys_0_instruction_master_translator:av_readdata -> nios2_qsys_0:i_readdata
	wire          nios2_qsys_0_instruction_master_readdatavalid;                                                                                 // nios2_qsys_0_instruction_master_translator:av_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire          nios2_qsys_0_data_master_waitrequest;                                                                                          // nios2_qsys_0_data_master_translator:av_waitrequest -> nios2_qsys_0:d_waitrequest
	wire   [31:0] nios2_qsys_0_data_master_writedata;                                                                                            // nios2_qsys_0:d_writedata -> nios2_qsys_0_data_master_translator:av_writedata
	wire   [26:0] nios2_qsys_0_data_master_address;                                                                                              // nios2_qsys_0:d_address -> nios2_qsys_0_data_master_translator:av_address
	wire          nios2_qsys_0_data_master_write;                                                                                                // nios2_qsys_0:d_write -> nios2_qsys_0_data_master_translator:av_write
	wire          nios2_qsys_0_data_master_read;                                                                                                 // nios2_qsys_0:d_read -> nios2_qsys_0_data_master_translator:av_read
	wire   [31:0] nios2_qsys_0_data_master_readdata;                                                                                             // nios2_qsys_0_data_master_translator:av_readdata -> nios2_qsys_0:d_readdata
	wire          nios2_qsys_0_data_master_debugaccess;                                                                                          // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_0_data_master_translator:av_debugaccess
	wire          nios2_qsys_0_data_master_readdatavalid;                                                                                        // nios2_qsys_0_data_master_translator:av_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire    [3:0] nios2_qsys_0_data_master_byteenable;                                                                                           // nios2_qsys_0:d_byteenable -> nios2_qsys_0_data_master_translator:av_byteenable
	wire          amd_0_avalon_master_waitrequest;                                                                                               // amd_0_avalon_master_translator:av_waitrequest -> amd_0:master_waitreq
	wire   [31:0] amd_0_avalon_master_address;                                                                                                   // amd_0:master_addr -> amd_0_avalon_master_translator:av_address
	wire   [15:0] amd_0_avalon_master_writedata;                                                                                                 // amd_0:master_wrdata -> amd_0_avalon_master_translator:av_writedata
	wire          amd_0_avalon_master_write;                                                                                                     // amd_0:master_write -> amd_0_avalon_master_translator:av_write
	wire          amd_0_avalon_master_read;                                                                                                      // amd_0:master_read -> amd_0_avalon_master_translator:av_read
	wire   [15:0] amd_0_avalon_master_readdata;                                                                                                  // amd_0_avalon_master_translator:av_readdata -> amd_0:master_rdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                                     // nios2_qsys_0:jtag_debug_module_waitrequest -> nios2_qsys_0_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                                       // nios2_qsys_0_jtag_debug_module_translator:av_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire    [8:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address;                                                         // nios2_qsys_0_jtag_debug_module_translator:av_address -> nios2_qsys_0:jtag_debug_module_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write;                                                           // nios2_qsys_0_jtag_debug_module_translator:av_write -> nios2_qsys_0:jtag_debug_module_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read;                                                            // nios2_qsys_0_jtag_debug_module_translator:av_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                                        // nios2_qsys_0:jtag_debug_module_readdata -> nios2_qsys_0_jtag_debug_module_translator:av_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                                     // nios2_qsys_0_jtag_debug_module_translator:av_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                                      // nios2_qsys_0_jtag_debug_module_translator:av_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire          new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest;                                                          // new_sdram_controller_0:za_waitrequest -> new_sdram_controller_0_s1_translator:av_waitrequest
	wire   [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata;                                                            // new_sdram_controller_0_s1_translator:av_writedata -> new_sdram_controller_0:az_data
	wire   [21:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address;                                                              // new_sdram_controller_0_s1_translator:av_address -> new_sdram_controller_0:az_addr
	wire          new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect;                                                           // new_sdram_controller_0_s1_translator:av_chipselect -> new_sdram_controller_0:az_cs
	wire          new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write;                                                                // new_sdram_controller_0_s1_translator:av_write -> new_sdram_controller_0:az_wr_n
	wire          new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read;                                                                 // new_sdram_controller_0_s1_translator:av_read -> new_sdram_controller_0:az_rd_n
	wire   [15:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata;                                                             // new_sdram_controller_0:za_data -> new_sdram_controller_0_s1_translator:av_readdata
	wire          new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid;                                                        // new_sdram_controller_0:za_valid -> new_sdram_controller_0_s1_translator:av_readdatavalid
	wire    [1:0] new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable;                                                           // new_sdram_controller_0_s1_translator:av_byteenable -> new_sdram_controller_0:az_be_n
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata;                                                                  // onchip_memory2_0_s1_translator:av_writedata -> onchip_memory2_0:writedata
	wire    [9:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_address;                                                                    // onchip_memory2_0_s1_translator:av_address -> onchip_memory2_0:address
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect;                                                                 // onchip_memory2_0_s1_translator:av_chipselect -> onchip_memory2_0:chipselect
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken;                                                                      // onchip_memory2_0_s1_translator:av_clken -> onchip_memory2_0:clken
	wire          onchip_memory2_0_s1_translator_avalon_anti_slave_0_write;                                                                      // onchip_memory2_0_s1_translator:av_write -> onchip_memory2_0:write
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata;                                                                   // onchip_memory2_0:readdata -> onchip_memory2_0_s1_translator:av_readdata
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable;                                                                 // onchip_memory2_0_s1_translator:av_byteenable -> onchip_memory2_0:byteenable
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest;                                              // to_external_bus_bridge_0:avalon_waitrequest -> to_external_bus_bridge_0_avalon_slave_translator:av_waitrequest
	wire   [15:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_writedata;                                                // to_external_bus_bridge_0_avalon_slave_translator:av_writedata -> to_external_bus_bridge_0:avalon_writedata
	wire   [14:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_address;                                                  // to_external_bus_bridge_0_avalon_slave_translator:av_address -> to_external_bus_bridge_0:avalon_address
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_chipselect;                                               // to_external_bus_bridge_0_avalon_slave_translator:av_chipselect -> to_external_bus_bridge_0:avalon_chipselect
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_write;                                                    // to_external_bus_bridge_0_avalon_slave_translator:av_write -> to_external_bus_bridge_0:avalon_write
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_read;                                                     // to_external_bus_bridge_0_avalon_slave_translator:av_read -> to_external_bus_bridge_0:avalon_read
	wire   [15:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_readdata;                                                 // to_external_bus_bridge_0:avalon_readdata -> to_external_bus_bridge_0_avalon_slave_translator:av_readdata
	wire    [1:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_byteenable;                                               // to_external_bus_bridge_0_avalon_slave_translator:av_byteenable -> to_external_bus_bridge_0:avalon_byteenable
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata;                                                           // rs232_0_avalon_rs232_slave_translator:av_writedata -> rs232_0:writedata
	wire    [0:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address;                                                             // rs232_0_avalon_rs232_slave_translator:av_address -> rs232_0:address
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect;                                                          // rs232_0_avalon_rs232_slave_translator:av_chipselect -> rs232_0:chipselect
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write;                                                               // rs232_0_avalon_rs232_slave_translator:av_write -> rs232_0:write
	wire          rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read;                                                                // rs232_0_avalon_rs232_slave_translator:av_read -> rs232_0:read
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata;                                                            // rs232_0:readdata -> rs232_0_avalon_rs232_slave_translator:av_readdata
	wire    [3:0] rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable;                                                          // rs232_0_avalon_rs232_slave_translator:av_byteenable -> rs232_0:byteenable
	wire    [1:0] pio_0_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_0_s1_translator:av_address -> pio_0:address
	wire   [31:0] pio_0_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_0:readdata -> pio_0_s1_translator:av_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest;                                                   // character_lcd_0:waitrequest -> character_lcd_0_avalon_lcd_slave_translator:av_waitrequest
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata;                                                     // character_lcd_0_avalon_lcd_slave_translator:av_writedata -> character_lcd_0:writedata
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address;                                                       // character_lcd_0_avalon_lcd_slave_translator:av_address -> character_lcd_0:address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect;                                                    // character_lcd_0_avalon_lcd_slave_translator:av_chipselect -> character_lcd_0:chipselect
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write;                                                         // character_lcd_0_avalon_lcd_slave_translator:av_write -> character_lcd_0:write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read;                                                          // character_lcd_0_avalon_lcd_slave_translator:av_read -> character_lcd_0:read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata;                                                      // character_lcd_0:readdata -> character_lcd_0_avalon_lcd_slave_translator:av_readdata
	wire    [1:0] pio_3_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_3_s1_translator:av_address -> pio_3:address
	wire   [31:0] pio_3_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_3:readdata -> pio_3_s1_translator:av_readdata
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                                                           // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire    [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                                             // timer_0_s1_translator:av_address -> timer_0:address
	wire          timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                                                          // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire          timer_0_s1_translator_avalon_anti_slave_0_write;                                                                               // timer_0_s1_translator:av_write -> timer_0:write_n
	wire   [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                                            // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_writedata;                                                                           // timer_1_s1_translator:av_writedata -> timer_1:writedata
	wire    [2:0] timer_1_s1_translator_avalon_anti_slave_0_address;                                                                             // timer_1_s1_translator:av_address -> timer_1:address
	wire          timer_1_s1_translator_avalon_anti_slave_0_chipselect;                                                                          // timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	wire          timer_1_s1_translator_avalon_anti_slave_0_write;                                                                               // timer_1_s1_translator:av_write -> timer_1:write_n
	wire   [15:0] timer_1_s1_translator_avalon_anti_slave_0_readdata;                                                                            // timer_1:readdata -> timer_1_s1_translator:av_readdata
	wire   [31:0] pio_4_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_4_s1_translator:av_writedata -> pio_4:writedata
	wire    [1:0] pio_4_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_4_s1_translator:av_address -> pio_4:address
	wire          pio_4_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_4_s1_translator:av_chipselect -> pio_4:chipselect
	wire          pio_4_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_4_s1_translator:av_write -> pio_4:write_n
	wire   [31:0] pio_4_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_4:readdata -> pio_4_s1_translator:av_readdata
	wire   [31:0] pio_5_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_5_s1_translator:av_writedata -> pio_5:writedata
	wire    [1:0] pio_5_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_5_s1_translator:av_address -> pio_5:address
	wire          pio_5_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_5_s1_translator:av_chipselect -> pio_5:chipselect
	wire          pio_5_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_5_s1_translator:av_write -> pio_5:write_n
	wire   [31:0] pio_5_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_5:readdata -> pio_5_s1_translator:av_readdata
	wire   [31:0] pio_6_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_6_s1_translator:av_writedata -> pio_6:writedata
	wire    [1:0] pio_6_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_6_s1_translator:av_address -> pio_6:address
	wire          pio_6_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_6_s1_translator:av_chipselect -> pio_6:chipselect
	wire          pio_6_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_6_s1_translator:av_write -> pio_6:write_n
	wire   [31:0] pio_6_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_6:readdata -> pio_6_s1_translator:av_readdata
	wire   [31:0] pio_7_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_7_s1_translator:av_writedata -> pio_7:writedata
	wire    [1:0] pio_7_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_7_s1_translator:av_address -> pio_7:address
	wire          pio_7_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_7_s1_translator:av_chipselect -> pio_7:chipselect
	wire          pio_7_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_7_s1_translator:av_write -> pio_7:write_n
	wire   [31:0] pio_7_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_7:readdata -> pio_7_s1_translator:av_readdata
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest;                           // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_waitrequest
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata;                             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_writedata -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_writedata
	wire    [7:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address;                               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_address -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_address
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect;                            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_chipselect -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_chip_select
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write;                                 // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_write -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_write
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read;                                  // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_read -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_read
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata;                              // Altera_UP_SD_Card_Avalon_Interface_0:o_avalon_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_readdata
	wire    [3:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable;                            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:av_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0:i_avalon_byteenable
	wire   [15:0] amd_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                                                                 // amd_0_avalon_slave_0_translator:av_writedata -> amd_0:slv_data
	wire   [15:0] amd_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                                                                   // amd_0_avalon_slave_0_translator:av_address -> amd_0:slv_addr
	wire          amd_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                                                     // amd_0_avalon_slave_0_translator:av_write -> amd_0:slv_start
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                                      // jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                                        // jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	wire    [0:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                                          // jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                                       // jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                                            // jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0:av_write_n
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                                             // jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0:av_read_n
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                                         // jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] pio_1_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_1_s1_translator:av_writedata -> pio_1:writedata
	wire    [1:0] pio_1_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_1_s1_translator:av_address -> pio_1:address
	wire          pio_1_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_1_s1_translator:av_chipselect -> pio_1:chipselect
	wire          pio_1_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_1_s1_translator:av_write -> pio_1:write_n
	wire   [31:0] pio_1_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_1:readdata -> pio_1_s1_translator:av_readdata
	wire   [31:0] pio_2_s1_translator_avalon_anti_slave_0_writedata;                                                                             // pio_2_s1_translator:av_writedata -> pio_2:writedata
	wire    [1:0] pio_2_s1_translator_avalon_anti_slave_0_address;                                                                               // pio_2_s1_translator:av_address -> pio_2:address
	wire          pio_2_s1_translator_avalon_anti_slave_0_chipselect;                                                                            // pio_2_s1_translator:av_chipselect -> pio_2:chipselect
	wire          pio_2_s1_translator_avalon_anti_slave_0_write;                                                                                 // pio_2_s1_translator:av_write -> pio_2:write_n
	wire   [31:0] pio_2_s1_translator_avalon_anti_slave_0_readdata;                                                                              // pio_2:readdata -> pio_2_s1_translator:av_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest;                                              // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_instruction_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount;                                               // nios2_qsys_0_instruction_master_translator:uav_burstcount -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata;                                                // nios2_qsys_0_instruction_master_translator:uav_writedata -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address;                                                  // nios2_qsys_0_instruction_master_translator:uav_address -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock;                                                     // nios2_qsys_0_instruction_master_translator:uav_lock -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write;                                                    // nios2_qsys_0_instruction_master_translator:uav_write -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read;                                                     // nios2_qsys_0_instruction_master_translator:uav_read -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata;                                                 // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_instruction_master_translator:uav_readdata
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess;                                              // nios2_qsys_0_instruction_master_translator:uav_debugaccess -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable;                                               // nios2_qsys_0_instruction_master_translator:uav_byteenable -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid;                                            // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_instruction_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest;                                                     // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_0_data_master_translator:uav_waitrequest
	wire    [2:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount;                                                      // nios2_qsys_0_data_master_translator:uav_burstcount -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata;                                                       // nios2_qsys_0_data_master_translator:uav_writedata -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_address;                                                         // nios2_qsys_0_data_master_translator:uav_address -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock;                                                            // nios2_qsys_0_data_master_translator:uav_lock -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_write;                                                           // nios2_qsys_0_data_master_translator:uav_write -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_read;                                                            // nios2_qsys_0_data_master_translator:uav_read -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata;                                                        // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_0_data_master_translator:uav_readdata
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess;                                                     // nios2_qsys_0_data_master_translator:uav_debugaccess -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable;                                                      // nios2_qsys_0_data_master_translator:uav_byteenable -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid;                                                   // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_0_data_master_translator:uav_readdatavalid
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                                                          // amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> amd_0_avalon_master_translator:uav_waitrequest
	wire    [1:0] amd_0_avalon_master_translator_avalon_universal_master_0_burstcount;                                                           // amd_0_avalon_master_translator:uav_burstcount -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [15:0] amd_0_avalon_master_translator_avalon_universal_master_0_writedata;                                                            // amd_0_avalon_master_translator:uav_writedata -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] amd_0_avalon_master_translator_avalon_universal_master_0_address;                                                              // amd_0_avalon_master_translator:uav_address -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_lock;                                                                 // amd_0_avalon_master_translator:uav_lock -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_write;                                                                // amd_0_avalon_master_translator:uav_write -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_read;                                                                 // amd_0_avalon_master_translator:uav_read -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [15:0] amd_0_avalon_master_translator_avalon_universal_master_0_readdata;                                                             // amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> amd_0_avalon_master_translator:uav_readdata
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                                                          // amd_0_avalon_master_translator:uav_debugaccess -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [1:0] amd_0_avalon_master_translator_avalon_universal_master_0_byteenable;                                                           // amd_0_avalon_master_translator:uav_byteenable -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                                                        // amd_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> amd_0_avalon_master_translator:uav_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                       // nios2_qsys_0_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_0_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                                         // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_0_jtag_debug_module_translator:uav_writedata
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_0_jtag_debug_module_translator:uav_address
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                                             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_0_jtag_debug_module_translator:uav_write
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_0_jtag_debug_module_translator:uav_lock
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_0_jtag_debug_module_translator:uav_read
	wire   [31:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                                          // nios2_qsys_0_jtag_debug_module_translator:uav_readdata -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                     // nios2_qsys_0_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_0_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_0_jtag_debug_module_translator:uav_byteenable
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                                      // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                           // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                    // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                   // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                  // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                 // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                            // new_sdram_controller_0_s1_translator:uav_waitrequest -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> new_sdram_controller_0_s1_translator:uav_burstcount
	wire   [15:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                              // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> new_sdram_controller_0_s1_translator:uav_writedata
	wire   [31:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> new_sdram_controller_0_s1_translator:uav_address
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                  // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> new_sdram_controller_0_s1_translator:uav_write
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> new_sdram_controller_0_s1_translator:uav_lock
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> new_sdram_controller_0_s1_translator:uav_read
	wire   [15:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                               // new_sdram_controller_0_s1_translator:uav_readdata -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                          // new_sdram_controller_0_s1_translator:uav_readdatavalid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> new_sdram_controller_0_s1_translator:uav_debugaccess
	wire    [1:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                             // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> new_sdram_controller_0_s1_translator:uav_byteenable
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                     // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                           // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                           // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                  // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                        // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                         // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                        // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                                      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                                       // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                                      // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                  // onchip_memory2_0_s1_translator:uav_waitrequest -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory2_0_s1_translator:uav_burstcount
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory2_0_s1_translator:uav_writedata
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory2_0_s1_translator:uav_address
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory2_0_s1_translator:uav_write
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory2_0_s1_translator:uav_lock
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory2_0_s1_translator:uav_read
	wire   [31:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                     // onchip_memory2_0_s1_translator:uav_readdata -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                // onchip_memory2_0_s1_translator:uav_readdatavalid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory2_0_s1_translator:uav_debugaccess
	wire    [3:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                   // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory2_0_s1_translator:uav_byteenable
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                           // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                 // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                      // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                               // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                              // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                             // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                            // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // to_external_bus_bridge_0_avalon_slave_translator:uav_waitrequest -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> to_external_bus_bridge_0_avalon_slave_translator:uav_burstcount
	wire   [15:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> to_external_bus_bridge_0_avalon_slave_translator:uav_writedata
	wire   [31:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                                    // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> to_external_bus_bridge_0_avalon_slave_translator:uav_address
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                                      // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> to_external_bus_bridge_0_avalon_slave_translator:uav_write
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                       // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> to_external_bus_bridge_0_avalon_slave_translator:uav_lock
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                                       // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> to_external_bus_bridge_0_avalon_slave_translator:uav_read
	wire   [15:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // to_external_bus_bridge_0_avalon_slave_translator:uav_readdata -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // to_external_bus_bridge_0_avalon_slave_translator:uav_readdatavalid -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> to_external_bus_bridge_0_avalon_slave_translator:uav_debugaccess
	wire    [1:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> to_external_bus_bridge_0_avalon_slave_translator:uav_byteenable
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                           // rs232_0_avalon_rs232_slave_translator:uav_waitrequest -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                            // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> rs232_0_avalon_rs232_slave_translator:uav_burstcount
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                             // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> rs232_0_avalon_rs232_slave_translator:uav_writedata
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address;                                               // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_address -> rs232_0_avalon_rs232_slave_translator:uav_address
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write;                                                 // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_write -> rs232_0_avalon_rs232_slave_translator:uav_write
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                                  // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_lock -> rs232_0_avalon_rs232_slave_translator:uav_lock
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read;                                                  // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_read -> rs232_0_avalon_rs232_slave_translator:uav_read
	wire   [31:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                              // rs232_0_avalon_rs232_slave_translator:uav_readdata -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                         // rs232_0_avalon_rs232_slave_translator:uav_readdatavalid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                           // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> rs232_0_avalon_rs232_slave_translator:uav_debugaccess
	wire    [3:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                            // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> rs232_0_avalon_rs232_slave_translator:uav_byteenable
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                    // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                          // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                  // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                           // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                          // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                 // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                       // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                               // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                        // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                       // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                     // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                      // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                     // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_0_s1_translator:uav_waitrequest -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_0_s1_translator:uav_burstcount
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_0_s1_translator:uav_writedata
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_0_s1_translator:uav_address
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_0_s1_translator:uav_write
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_0_s1_translator:uav_lock
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_0_s1_translator:uav_read
	wire   [31:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_0_s1_translator:uav_readdata -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_0_s1_translator:uav_readdatavalid -> pio_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_0_s1_translator:uav_debugaccess
	wire    [3:0] pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_0_s1_translator:uav_byteenable
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // character_lcd_0_avalon_lcd_slave_translator:uav_waitrequest -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> character_lcd_0_avalon_lcd_slave_translator:uav_burstcount
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> character_lcd_0_avalon_lcd_slave_translator:uav_writedata
	wire   [31:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address;                                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_address -> character_lcd_0_avalon_lcd_slave_translator:uav_address
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write;                                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_write -> character_lcd_0_avalon_lcd_slave_translator:uav_write
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_lock -> character_lcd_0_avalon_lcd_slave_translator:uav_lock
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read;                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_read -> character_lcd_0_avalon_lcd_slave_translator:uav_read
	wire    [7:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // character_lcd_0_avalon_lcd_slave_translator:uav_readdata -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // character_lcd_0_avalon_lcd_slave_translator:uav_readdatavalid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> character_lcd_0_avalon_lcd_slave_translator:uav_debugaccess
	wire    [0:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> character_lcd_0_avalon_lcd_slave_translator:uav_byteenable
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [82:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [82:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire    [9:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_3_s1_translator:uav_waitrequest -> pio_3_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_3_s1_translator:uav_burstcount
	wire   [31:0] pio_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_3_s1_translator:uav_writedata
	wire   [31:0] pio_3_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_3_s1_translator:uav_address
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_3_s1_translator:uav_write
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_3_s1_translator:uav_lock
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_3_s1_translator:uav_read
	wire   [31:0] pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_3_s1_translator:uav_readdata -> pio_3_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_3_s1_translator:uav_readdatavalid -> pio_3_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_3_s1_translator:uav_debugaccess
	wire    [3:0] pio_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_3_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_3_s1_translator:uav_byteenable
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_3_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_3_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_3_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_3_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_3_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_3_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_3_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                           // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                            // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                             // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                               // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire   [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                              // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                         // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire    [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                            // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                          // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                 // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                       // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                               // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                        // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                       // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                           // timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                            // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                             // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                               // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	wire   [31:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                              // timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                         // timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	wire    [3:0] timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                            // timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                          // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                          // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                 // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                       // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                               // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                        // timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                       // timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                      // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                     // timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_4_s1_translator:uav_waitrequest -> pio_4_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_4_s1_translator:uav_burstcount
	wire   [31:0] pio_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_4_s1_translator:uav_writedata
	wire   [31:0] pio_4_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_4_s1_translator:uav_address
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_4_s1_translator:uav_write
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_4_s1_translator:uav_lock
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_4_s1_translator:uav_read
	wire   [31:0] pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_4_s1_translator:uav_readdata -> pio_4_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_4_s1_translator:uav_readdatavalid -> pio_4_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_4_s1_translator:uav_debugaccess
	wire    [3:0] pio_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_4_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_4_s1_translator:uav_byteenable
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_4_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_4_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_4_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_4_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_4_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_4_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_4_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_5_s1_translator:uav_waitrequest -> pio_5_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_5_s1_translator:uav_burstcount
	wire   [31:0] pio_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_5_s1_translator:uav_writedata
	wire   [31:0] pio_5_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_5_s1_translator:uav_address
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_5_s1_translator:uav_write
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_5_s1_translator:uav_lock
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_5_s1_translator:uav_read
	wire   [31:0] pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_5_s1_translator:uav_readdata -> pio_5_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_5_s1_translator:uav_readdatavalid -> pio_5_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_5_s1_translator:uav_debugaccess
	wire    [3:0] pio_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_5_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_5_s1_translator:uav_byteenable
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_5_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_5_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_5_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_5_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_5_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_5_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_5_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_6_s1_translator:uav_waitrequest -> pio_6_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_6_s1_translator:uav_burstcount
	wire   [31:0] pio_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_6_s1_translator:uav_writedata
	wire   [31:0] pio_6_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_6_s1_translator:uav_address
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_6_s1_translator:uav_write
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_6_s1_translator:uav_lock
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_6_s1_translator:uav_read
	wire   [31:0] pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_6_s1_translator:uav_readdata -> pio_6_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_6_s1_translator:uav_readdatavalid -> pio_6_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_6_s1_translator:uav_debugaccess
	wire    [3:0] pio_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_6_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_6_s1_translator:uav_byteenable
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_6_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_6_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_6_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_6_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_6_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_6_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_6_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_7_s1_translator:uav_waitrequest -> pio_7_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_7_s1_translator:uav_burstcount
	wire   [31:0] pio_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_7_s1_translator:uav_writedata
	wire   [31:0] pio_7_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_7_s1_translator:uav_address
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_7_s1_translator:uav_write
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_7_s1_translator:uav_lock
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_7_s1_translator:uav_read
	wire   [31:0] pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_7_s1_translator:uav_readdata -> pio_7_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_7_s1_translator:uav_readdatavalid -> pio_7_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_7_s1_translator:uav_debugaccess
	wire    [3:0] pio_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_7_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_7_s1_translator:uav_byteenable
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_7_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_7_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_7_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_7_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_7_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_7_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_7_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_waitrequest -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_burstcount
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_writedata
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_address -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_address
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_write -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_write
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_lock -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_lock
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_read -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_read
	wire   [31:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdata -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_readdatavalid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_debugaccess
	wire    [3:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:uav_byteenable
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                 // amd_0_avalon_slave_0_translator:uav_waitrequest -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                  // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> amd_0_avalon_slave_0_translator:uav_burstcount
	wire   [15:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;                                                   // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> amd_0_avalon_slave_0_translator:uav_writedata
	wire   [31:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                                                     // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> amd_0_avalon_slave_0_translator:uav_address
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                                                       // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> amd_0_avalon_slave_0_translator:uav_write
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                                                        // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> amd_0_avalon_slave_0_translator:uav_lock
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                                                        // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> amd_0_avalon_slave_0_translator:uav_read
	wire   [15:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                                                    // amd_0_avalon_slave_0_translator:uav_readdata -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                               // amd_0_avalon_slave_0_translator:uav_readdatavalid -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                 // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> amd_0_avalon_slave_0_translator:uav_debugaccess
	wire    [1:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                  // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> amd_0_avalon_slave_0_translator:uav_byteenable
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                          // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                        // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [91:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;                                                 // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                       // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                             // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                     // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [91:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                              // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                             // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                           // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                            // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                           // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                        // jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                          // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                           // jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                      // jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                         // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                 // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                       // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                            // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                     // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                    // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                   // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                  // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_1_s1_translator:uav_waitrequest -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_1_s1_translator:uav_burstcount
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_1_s1_translator:uav_writedata
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_1_s1_translator:uav_address
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_1_s1_translator:uav_write
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_1_s1_translator:uav_lock
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_1_s1_translator:uav_read
	wire   [31:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_1_s1_translator:uav_readdata -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_1_s1_translator:uav_readdatavalid -> pio_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_1_s1_translator:uav_debugaccess
	wire    [3:0] pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_1_s1_translator:uav_byteenable
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                                             // pio_2_s1_translator:uav_waitrequest -> pio_2_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pio_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                                              // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_2_s1_translator:uav_burstcount
	wire   [31:0] pio_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                                               // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_2_s1_translator:uav_writedata
	wire   [31:0] pio_2_s1_translator_avalon_universal_slave_0_agent_m0_address;                                                                 // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_2_s1_translator:uav_address
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_write;                                                                   // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_2_s1_translator:uav_write
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                                                    // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_2_s1_translator:uav_lock
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_read;                                                                    // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_2_s1_translator:uav_read
	wire   [31:0] pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                                                // pio_2_s1_translator:uav_readdata -> pio_2_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                                           // pio_2_s1_translator:uav_readdatavalid -> pio_2_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                                             // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_2_s1_translator:uav_debugaccess
	wire    [3:0] pio_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                                              // pio_2_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_2_s1_translator:uav_byteenable
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                                                      // pio_2_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                                            // pio_2_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                                                    // pio_2_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [109:0] pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                                             // pio_2_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                                            // pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_2_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                                                   // pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                                         // pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                                                 // pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [109:0] pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                                          // pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                                         // pio_2_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                                                       // pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                                        // pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                                                       // pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_2_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                     // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                                           // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                   // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [108:0] nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                                            // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                                           // addr_router:sink_ready -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                            // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                                  // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                          // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [108:0] nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data;                                                   // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                                  // addr_router_001:sink_ready -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                                                 // amd_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                                                       // amd_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                                               // amd_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire   [90:0] amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                                                        // amd_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                                                       // addr_router_002:sink_ready -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                       // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                                             // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                     // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [108:0] nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                              // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                                             // id_router:sink_ready -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                            // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                  // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                          // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire   [90:0] new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                  // id_router_001:sink_ready -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                  // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                        // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [108:0] onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                         // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                        // id_router_002:sink_ready -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                      // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire   [90:0] to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                                       // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_003:sink_ready -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                           // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                                 // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                         // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [108:0] rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data;                                                  // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                                 // id_router_004:sink_ready -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [108:0] pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_005:sink_ready -> pio_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                           // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire   [81:0] character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data;                                            // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_006:sink_ready -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_3_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_3_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_3_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [108:0] pio_3_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_3_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          pio_3_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_007:sink_ready -> pio_3_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [108:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                  // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                 // id_router_008:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                           // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                 // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                         // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [108:0] timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                  // timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                 // id_router_009:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_4_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_4_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_4_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [108:0] pio_4_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_4_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          pio_4_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_010:sink_ready -> pio_4_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_5_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_5_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_5_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [108:0] pio_5_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_5_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          pio_5_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_011:sink_ready -> pio_5_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_6_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_6_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_6_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [108:0] pio_6_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_6_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          pio_6_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_012:sink_ready -> pio_6_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_7_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_7_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_7_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [108:0] pio_7_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_7_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pio_7_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_013:sink_ready -> pio_7_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire  [108:0] altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_014:sink_ready -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                 // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                                                       // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                               // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [90:0] amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                                                        // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                                                       // id_router_015:sink_ready -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                        // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                              // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                      // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire  [108:0] jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                                               // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                              // id_router_016:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire  [108:0] pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_017:sink_ready -> pio_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                                             // pio_2_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                                                   // pio_2_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                                           // pio_2_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire  [108:0] pio_2_s1_translator_avalon_universal_slave_0_agent_rp_data;                                                                    // pio_2_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          pio_2_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                                                   // id_router_018:sink_ready -> pio_2_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                                                   // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                                                         // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                                                 // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [108:0] addr_router_src_data;                                                                                                          // addr_router:src_data -> limiter:cmd_sink_data
	wire   [18:0] addr_router_src_channel;                                                                                                       // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                                                         // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                                                   // limiter:rsp_src_endofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                                         // limiter:rsp_src_valid -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                                                 // limiter:rsp_src_startofpacket -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] limiter_rsp_src_data;                                                                                                          // limiter:rsp_src_data -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_rsp_src_channel;                                                                                                       // limiter:rsp_src_channel -> nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                                         // nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                                               // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                                                     // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                                             // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [108:0] addr_router_001_src_data;                                                                                                      // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire   [18:0] addr_router_001_src_channel;                                                                                                   // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                                                     // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                                               // limiter_001:rsp_src_endofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                                                     // limiter_001:rsp_src_valid -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                                             // limiter_001:rsp_src_startofpacket -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [108:0] limiter_001_rsp_src_data;                                                                                                      // limiter_001:rsp_src_data -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] limiter_001_rsp_src_channel;                                                                                                   // limiter_001:rsp_src_channel -> nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                                                     // nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                                             // burst_adapter:source0_endofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                                                   // burst_adapter:source0_valid -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                                           // burst_adapter:source0_startofpacket -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_source0_data;                                                                                                    // burst_adapter:source0_data -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                                                   // new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire   [18:0] burst_adapter_source0_channel;                                                                                                 // burst_adapter:source0_channel -> new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                                                         // burst_adapter_001:source0_endofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                                               // burst_adapter_001:source0_valid -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                                                       // burst_adapter_001:source0_startofpacket -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_001_source0_data;                                                                                                // burst_adapter_001:source0_data -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                                               // to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire   [18:0] burst_adapter_001_source0_channel;                                                                                             // burst_adapter_001:source0_channel -> to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                                                         // burst_adapter_002:source0_endofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                                               // burst_adapter_002:source0_valid -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                                                       // burst_adapter_002:source0_startofpacket -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [81:0] burst_adapter_002_source0_data;                                                                                                // burst_adapter_002:source0_data -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                                               // character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire   [18:0] burst_adapter_002_source0_channel;                                                                                             // burst_adapter_002:source0_channel -> character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                                                         // burst_adapter_003:source0_endofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                                               // burst_adapter_003:source0_valid -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                                                       // burst_adapter_003:source0_startofpacket -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [90:0] burst_adapter_003_source0_data;                                                                                                // burst_adapter_003:source0_data -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                                               // amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire   [18:0] burst_adapter_003_source0_channel;                                                                                             // burst_adapter_003:source0_channel -> amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                                                // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, character_lcd_0:reset, character_lcd_0_avalon_lcd_slave_translator:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent:reset, character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, cmd_xbar_mux_009:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, irq_mapper:reset, jtag_uart_0:rst_n, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, new_sdram_controller_0:reset_n, new_sdram_controller_0_s1_translator:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, nios2_qsys_0:reset_n, nios2_qsys_0_data_master_translator:reset, nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_instruction_master_translator:reset, nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory2_0:reset, onchip_memory2_0_s1_translator:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_0:reset_n, pio_0_s1_translator:reset, pio_0_s1_translator_avalon_universal_slave_0_agent:reset, pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_1:reset_n, pio_1_s1_translator:reset, pio_1_s1_translator_avalon_universal_slave_0_agent:reset, pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_2:reset_n, pio_2_s1_translator:reset, pio_2_s1_translator_avalon_universal_slave_0_agent:reset, pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_3:reset_n, pio_3_s1_translator:reset, pio_3_s1_translator_avalon_universal_slave_0_agent:reset, pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rs232_0:reset, rs232_0_avalon_rs232_slave_translator:reset, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:reset, rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1:reset_n, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, to_external_bus_bridge_0:reset, to_external_bus_bridge_0_avalon_slave_translator:reset, to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset, width_adapter_012:reset, width_adapter_013:reset]
	wire          rst_controller_reset_out_reset_req;                                                                                            // rst_controller:reset_req -> onchip_memory2_0:reset_req
	wire          nios2_qsys_0_jtag_debug_module_reset_reset;                                                                                    // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                                                                            // rst_controller_001:reset_out -> up_clocks_0:reset
	wire          rst_controller_002_reset_out_reset;                                                                                            // rst_controller_002:reset_out -> [Altera_UP_SD_Card_Avalon_Interface_0:i_reset_n, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:reset, Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router_002:reset, amd_0:reset_n, amd_0_avalon_master_translator:reset, amd_0_avalon_master_translator_avalon_universal_master_0_agent:reset, amd_0_avalon_slave_0_translator:reset, amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_003:reset, cmd_xbar_demux_002:reset, cmd_xbar_mux_010:reset, cmd_xbar_mux_011:reset, cmd_xbar_mux_012:reset, cmd_xbar_mux_013:reset, cmd_xbar_mux_014:reset, cmd_xbar_mux_015:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, pio_4:reset_n, pio_4_s1_translator:reset, pio_4_s1_translator_avalon_universal_slave_0_agent:reset, pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_5:reset_n, pio_5_s1_translator:reset, pio_5_s1_translator_avalon_universal_slave_0_agent:reset, pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_6:reset_n, pio_6_s1_translator:reset, pio_6_s1_translator_avalon_universal_slave_0_agent:reset, pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_7:reset_n, pio_7_s1_translator:reset, pio_7_s1_translator_avalon_universal_slave_0_agent:reset, pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux_002:reset, width_adapter_014:reset, width_adapter_015:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                                               // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                                                     // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                                             // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src0_data;                                                                                                      // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire   [18:0] cmd_xbar_demux_src0_channel;                                                                                                   // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire          cmd_xbar_demux_src0_ready;                                                                                                     // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src2_endofpacket;                                                                                               // cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                                                                     // cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                                                             // cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src2_data;                                                                                                      // cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	wire   [18:0] cmd_xbar_demux_src2_channel;                                                                                                   // cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_src2_ready;                                                                                                     // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	wire          cmd_xbar_demux_src4_endofpacket;                                                                                               // cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_src4_valid;                                                                                                     // cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_src4_startofpacket;                                                                                             // cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src4_data;                                                                                                      // cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	wire   [18:0] cmd_xbar_demux_src4_channel;                                                                                                   // cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_src4_ready;                                                                                                     // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	wire          cmd_xbar_demux_src5_endofpacket;                                                                                               // cmd_xbar_demux:src5_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_src5_valid;                                                                                                     // cmd_xbar_demux:src5_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_src5_startofpacket;                                                                                             // cmd_xbar_demux:src5_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src5_data;                                                                                                      // cmd_xbar_demux:src5_data -> cmd_xbar_mux_005:sink0_data
	wire   [18:0] cmd_xbar_demux_src5_channel;                                                                                                   // cmd_xbar_demux:src5_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_src5_ready;                                                                                                     // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux:src5_ready
	wire          cmd_xbar_demux_src7_endofpacket;                                                                                               // cmd_xbar_demux:src7_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire          cmd_xbar_demux_src7_valid;                                                                                                     // cmd_xbar_demux:src7_valid -> cmd_xbar_mux_007:sink0_valid
	wire          cmd_xbar_demux_src7_startofpacket;                                                                                             // cmd_xbar_demux:src7_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src7_data;                                                                                                      // cmd_xbar_demux:src7_data -> cmd_xbar_mux_007:sink0_data
	wire   [18:0] cmd_xbar_demux_src7_channel;                                                                                                   // cmd_xbar_demux:src7_channel -> cmd_xbar_mux_007:sink0_channel
	wire          cmd_xbar_demux_src7_ready;                                                                                                     // cmd_xbar_mux_007:sink0_ready -> cmd_xbar_demux:src7_ready
	wire          cmd_xbar_demux_src8_endofpacket;                                                                                               // cmd_xbar_demux:src8_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          cmd_xbar_demux_src8_valid;                                                                                                     // cmd_xbar_demux:src8_valid -> cmd_xbar_mux_008:sink0_valid
	wire          cmd_xbar_demux_src8_startofpacket;                                                                                             // cmd_xbar_demux:src8_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src8_data;                                                                                                      // cmd_xbar_demux:src8_data -> cmd_xbar_mux_008:sink0_data
	wire   [18:0] cmd_xbar_demux_src8_channel;                                                                                                   // cmd_xbar_demux:src8_channel -> cmd_xbar_mux_008:sink0_channel
	wire          cmd_xbar_demux_src8_ready;                                                                                                     // cmd_xbar_mux_008:sink0_ready -> cmd_xbar_demux:src8_ready
	wire          cmd_xbar_demux_src9_endofpacket;                                                                                               // cmd_xbar_demux:src9_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          cmd_xbar_demux_src9_valid;                                                                                                     // cmd_xbar_demux:src9_valid -> cmd_xbar_mux_009:sink0_valid
	wire          cmd_xbar_demux_src9_startofpacket;                                                                                             // cmd_xbar_demux:src9_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src9_data;                                                                                                      // cmd_xbar_demux:src9_data -> cmd_xbar_mux_009:sink0_data
	wire   [18:0] cmd_xbar_demux_src9_channel;                                                                                                   // cmd_xbar_demux:src9_channel -> cmd_xbar_mux_009:sink0_channel
	wire          cmd_xbar_demux_src9_ready;                                                                                                     // cmd_xbar_mux_009:sink0_ready -> cmd_xbar_demux:src9_ready
	wire          cmd_xbar_demux_src10_endofpacket;                                                                                              // cmd_xbar_demux:src10_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          cmd_xbar_demux_src10_valid;                                                                                                    // cmd_xbar_demux:src10_valid -> cmd_xbar_mux_010:sink0_valid
	wire          cmd_xbar_demux_src10_startofpacket;                                                                                            // cmd_xbar_demux:src10_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src10_data;                                                                                                     // cmd_xbar_demux:src10_data -> cmd_xbar_mux_010:sink0_data
	wire   [18:0] cmd_xbar_demux_src10_channel;                                                                                                  // cmd_xbar_demux:src10_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_src10_ready;                                                                                                    // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux:src10_ready
	wire          cmd_xbar_demux_src11_endofpacket;                                                                                              // cmd_xbar_demux:src11_endofpacket -> cmd_xbar_mux_011:sink0_endofpacket
	wire          cmd_xbar_demux_src11_valid;                                                                                                    // cmd_xbar_demux:src11_valid -> cmd_xbar_mux_011:sink0_valid
	wire          cmd_xbar_demux_src11_startofpacket;                                                                                            // cmd_xbar_demux:src11_startofpacket -> cmd_xbar_mux_011:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src11_data;                                                                                                     // cmd_xbar_demux:src11_data -> cmd_xbar_mux_011:sink0_data
	wire   [18:0] cmd_xbar_demux_src11_channel;                                                                                                  // cmd_xbar_demux:src11_channel -> cmd_xbar_mux_011:sink0_channel
	wire          cmd_xbar_demux_src11_ready;                                                                                                    // cmd_xbar_mux_011:sink0_ready -> cmd_xbar_demux:src11_ready
	wire          cmd_xbar_demux_src12_endofpacket;                                                                                              // cmd_xbar_demux:src12_endofpacket -> cmd_xbar_mux_012:sink0_endofpacket
	wire          cmd_xbar_demux_src12_valid;                                                                                                    // cmd_xbar_demux:src12_valid -> cmd_xbar_mux_012:sink0_valid
	wire          cmd_xbar_demux_src12_startofpacket;                                                                                            // cmd_xbar_demux:src12_startofpacket -> cmd_xbar_mux_012:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src12_data;                                                                                                     // cmd_xbar_demux:src12_data -> cmd_xbar_mux_012:sink0_data
	wire   [18:0] cmd_xbar_demux_src12_channel;                                                                                                  // cmd_xbar_demux:src12_channel -> cmd_xbar_mux_012:sink0_channel
	wire          cmd_xbar_demux_src12_ready;                                                                                                    // cmd_xbar_mux_012:sink0_ready -> cmd_xbar_demux:src12_ready
	wire          cmd_xbar_demux_src13_endofpacket;                                                                                              // cmd_xbar_demux:src13_endofpacket -> cmd_xbar_mux_013:sink0_endofpacket
	wire          cmd_xbar_demux_src13_valid;                                                                                                    // cmd_xbar_demux:src13_valid -> cmd_xbar_mux_013:sink0_valid
	wire          cmd_xbar_demux_src13_startofpacket;                                                                                            // cmd_xbar_demux:src13_startofpacket -> cmd_xbar_mux_013:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src13_data;                                                                                                     // cmd_xbar_demux:src13_data -> cmd_xbar_mux_013:sink0_data
	wire   [18:0] cmd_xbar_demux_src13_channel;                                                                                                  // cmd_xbar_demux:src13_channel -> cmd_xbar_mux_013:sink0_channel
	wire          cmd_xbar_demux_src13_ready;                                                                                                    // cmd_xbar_mux_013:sink0_ready -> cmd_xbar_demux:src13_ready
	wire          cmd_xbar_demux_src14_endofpacket;                                                                                              // cmd_xbar_demux:src14_endofpacket -> cmd_xbar_mux_014:sink0_endofpacket
	wire          cmd_xbar_demux_src14_valid;                                                                                                    // cmd_xbar_demux:src14_valid -> cmd_xbar_mux_014:sink0_valid
	wire          cmd_xbar_demux_src14_startofpacket;                                                                                            // cmd_xbar_demux:src14_startofpacket -> cmd_xbar_mux_014:sink0_startofpacket
	wire  [108:0] cmd_xbar_demux_src14_data;                                                                                                     // cmd_xbar_demux:src14_data -> cmd_xbar_mux_014:sink0_data
	wire   [18:0] cmd_xbar_demux_src14_channel;                                                                                                  // cmd_xbar_demux:src14_channel -> cmd_xbar_mux_014:sink0_channel
	wire          cmd_xbar_demux_src14_ready;                                                                                                    // cmd_xbar_mux_014:sink0_ready -> cmd_xbar_demux:src14_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                                           // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                                                 // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                                         // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src0_data;                                                                                                  // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src0_channel;                                                                                               // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                                                 // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                                           // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                                                 // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                                                         // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src2_data;                                                                                                  // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src2_channel;                                                                                               // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                                                 // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                                           // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                                                 // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                                                         // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src4_data;                                                                                                  // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src4_channel;                                                                                               // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                                                 // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                                           // cmd_xbar_demux_001:src5_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                                                 // cmd_xbar_demux_001:src5_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                                                         // cmd_xbar_demux_001:src5_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src5_data;                                                                                                  // cmd_xbar_demux_001:src5_data -> cmd_xbar_mux_005:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src5_channel;                                                                                               // cmd_xbar_demux_001:src5_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                                                 // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_001:src5_ready
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                                           // cmd_xbar_demux_001:src7_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                                                 // cmd_xbar_demux_001:src7_valid -> cmd_xbar_mux_007:sink1_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                                                         // cmd_xbar_demux_001:src7_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src7_data;                                                                                                  // cmd_xbar_demux_001:src7_data -> cmd_xbar_mux_007:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src7_channel;                                                                                               // cmd_xbar_demux_001:src7_channel -> cmd_xbar_mux_007:sink1_channel
	wire          cmd_xbar_demux_001_src7_ready;                                                                                                 // cmd_xbar_mux_007:sink1_ready -> cmd_xbar_demux_001:src7_ready
	wire          cmd_xbar_demux_001_src8_endofpacket;                                                                                           // cmd_xbar_demux_001:src8_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          cmd_xbar_demux_001_src8_valid;                                                                                                 // cmd_xbar_demux_001:src8_valid -> cmd_xbar_mux_008:sink1_valid
	wire          cmd_xbar_demux_001_src8_startofpacket;                                                                                         // cmd_xbar_demux_001:src8_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src8_data;                                                                                                  // cmd_xbar_demux_001:src8_data -> cmd_xbar_mux_008:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src8_channel;                                                                                               // cmd_xbar_demux_001:src8_channel -> cmd_xbar_mux_008:sink1_channel
	wire          cmd_xbar_demux_001_src8_ready;                                                                                                 // cmd_xbar_mux_008:sink1_ready -> cmd_xbar_demux_001:src8_ready
	wire          cmd_xbar_demux_001_src9_endofpacket;                                                                                           // cmd_xbar_demux_001:src9_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          cmd_xbar_demux_001_src9_valid;                                                                                                 // cmd_xbar_demux_001:src9_valid -> cmd_xbar_mux_009:sink1_valid
	wire          cmd_xbar_demux_001_src9_startofpacket;                                                                                         // cmd_xbar_demux_001:src9_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src9_data;                                                                                                  // cmd_xbar_demux_001:src9_data -> cmd_xbar_mux_009:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src9_channel;                                                                                               // cmd_xbar_demux_001:src9_channel -> cmd_xbar_mux_009:sink1_channel
	wire          cmd_xbar_demux_001_src9_ready;                                                                                                 // cmd_xbar_mux_009:sink1_ready -> cmd_xbar_demux_001:src9_ready
	wire          cmd_xbar_demux_001_src10_endofpacket;                                                                                          // cmd_xbar_demux_001:src10_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_001_src10_valid;                                                                                                // cmd_xbar_demux_001:src10_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_001_src10_startofpacket;                                                                                        // cmd_xbar_demux_001:src10_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src10_data;                                                                                                 // cmd_xbar_demux_001:src10_data -> cmd_xbar_mux_010:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src10_channel;                                                                                              // cmd_xbar_demux_001:src10_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_001_src10_ready;                                                                                                // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_001:src10_ready
	wire          cmd_xbar_demux_001_src11_endofpacket;                                                                                          // cmd_xbar_demux_001:src11_endofpacket -> cmd_xbar_mux_011:sink1_endofpacket
	wire          cmd_xbar_demux_001_src11_valid;                                                                                                // cmd_xbar_demux_001:src11_valid -> cmd_xbar_mux_011:sink1_valid
	wire          cmd_xbar_demux_001_src11_startofpacket;                                                                                        // cmd_xbar_demux_001:src11_startofpacket -> cmd_xbar_mux_011:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src11_data;                                                                                                 // cmd_xbar_demux_001:src11_data -> cmd_xbar_mux_011:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src11_channel;                                                                                              // cmd_xbar_demux_001:src11_channel -> cmd_xbar_mux_011:sink1_channel
	wire          cmd_xbar_demux_001_src11_ready;                                                                                                // cmd_xbar_mux_011:sink1_ready -> cmd_xbar_demux_001:src11_ready
	wire          cmd_xbar_demux_001_src12_endofpacket;                                                                                          // cmd_xbar_demux_001:src12_endofpacket -> cmd_xbar_mux_012:sink1_endofpacket
	wire          cmd_xbar_demux_001_src12_valid;                                                                                                // cmd_xbar_demux_001:src12_valid -> cmd_xbar_mux_012:sink1_valid
	wire          cmd_xbar_demux_001_src12_startofpacket;                                                                                        // cmd_xbar_demux_001:src12_startofpacket -> cmd_xbar_mux_012:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src12_data;                                                                                                 // cmd_xbar_demux_001:src12_data -> cmd_xbar_mux_012:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src12_channel;                                                                                              // cmd_xbar_demux_001:src12_channel -> cmd_xbar_mux_012:sink1_channel
	wire          cmd_xbar_demux_001_src12_ready;                                                                                                // cmd_xbar_mux_012:sink1_ready -> cmd_xbar_demux_001:src12_ready
	wire          cmd_xbar_demux_001_src13_endofpacket;                                                                                          // cmd_xbar_demux_001:src13_endofpacket -> cmd_xbar_mux_013:sink1_endofpacket
	wire          cmd_xbar_demux_001_src13_valid;                                                                                                // cmd_xbar_demux_001:src13_valid -> cmd_xbar_mux_013:sink1_valid
	wire          cmd_xbar_demux_001_src13_startofpacket;                                                                                        // cmd_xbar_demux_001:src13_startofpacket -> cmd_xbar_mux_013:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src13_data;                                                                                                 // cmd_xbar_demux_001:src13_data -> cmd_xbar_mux_013:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src13_channel;                                                                                              // cmd_xbar_demux_001:src13_channel -> cmd_xbar_mux_013:sink1_channel
	wire          cmd_xbar_demux_001_src13_ready;                                                                                                // cmd_xbar_mux_013:sink1_ready -> cmd_xbar_demux_001:src13_ready
	wire          cmd_xbar_demux_001_src14_endofpacket;                                                                                          // cmd_xbar_demux_001:src14_endofpacket -> cmd_xbar_mux_014:sink1_endofpacket
	wire          cmd_xbar_demux_001_src14_valid;                                                                                                // cmd_xbar_demux_001:src14_valid -> cmd_xbar_mux_014:sink1_valid
	wire          cmd_xbar_demux_001_src14_startofpacket;                                                                                        // cmd_xbar_demux_001:src14_startofpacket -> cmd_xbar_mux_014:sink1_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src14_data;                                                                                                 // cmd_xbar_demux_001:src14_data -> cmd_xbar_mux_014:sink1_data
	wire   [18:0] cmd_xbar_demux_001_src14_channel;                                                                                              // cmd_xbar_demux_001:src14_channel -> cmd_xbar_mux_014:sink1_channel
	wire          cmd_xbar_demux_001_src14_ready;                                                                                                // cmd_xbar_mux_014:sink1_ready -> cmd_xbar_demux_001:src14_ready
	wire          cmd_xbar_demux_001_src16_endofpacket;                                                                                          // cmd_xbar_demux_001:src16_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src16_valid;                                                                                                // cmd_xbar_demux_001:src16_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src16_startofpacket;                                                                                        // cmd_xbar_demux_001:src16_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src16_data;                                                                                                 // cmd_xbar_demux_001:src16_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src16_channel;                                                                                              // cmd_xbar_demux_001:src16_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src17_endofpacket;                                                                                          // cmd_xbar_demux_001:src17_endofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src17_valid;                                                                                                // cmd_xbar_demux_001:src17_valid -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src17_startofpacket;                                                                                        // cmd_xbar_demux_001:src17_startofpacket -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src17_data;                                                                                                 // cmd_xbar_demux_001:src17_data -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src17_channel;                                                                                              // cmd_xbar_demux_001:src17_channel -> pio_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_001_src18_endofpacket;                                                                                          // cmd_xbar_demux_001:src18_endofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_001_src18_valid;                                                                                                // cmd_xbar_demux_001:src18_valid -> pio_2_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_001_src18_startofpacket;                                                                                        // cmd_xbar_demux_001:src18_startofpacket -> pio_2_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src18_data;                                                                                                 // cmd_xbar_demux_001:src18_data -> pio_2_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_demux_001_src18_channel;                                                                                              // cmd_xbar_demux_001:src18_channel -> pio_2_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                                           // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                                                 // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                                         // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire   [90:0] cmd_xbar_demux_002_src0_data;                                                                                                  // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_001:sink2_data
	wire   [18:0] cmd_xbar_demux_002_src0_channel;                                                                                               // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                                                 // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                                           // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                                                 // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                                                         // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire   [90:0] cmd_xbar_demux_002_src1_data;                                                                                                  // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_003:sink2_data
	wire   [18:0] cmd_xbar_demux_002_src1_channel;                                                                                               // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                                                 // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_src0_endofpacket;                                                                                               // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                                                     // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                                             // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src0_data;                                                                                                      // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire   [18:0] rsp_xbar_demux_src0_channel;                                                                                                   // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                                                     // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                                               // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                                                     // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                                             // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [108:0] rsp_xbar_demux_src1_data;                                                                                                      // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire   [18:0] rsp_xbar_demux_src1_channel;                                                                                                   // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_src1_ready;                                                                                                     // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                                           // rsp_xbar_demux_001:src2_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                                                 // rsp_xbar_demux_001:src2_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                                         // rsp_xbar_demux_001:src2_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src2_data;                                                                                                  // rsp_xbar_demux_001:src2_data -> rsp_xbar_mux_002:sink0_data
	wire   [18:0] rsp_xbar_demux_001_src2_channel;                                                                                               // rsp_xbar_demux_001:src2_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                                                 // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                                           // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                                                 // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                                         // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [108:0] rsp_xbar_demux_002_src0_data;                                                                                                  // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire   [18:0] rsp_xbar_demux_002_src0_channel;                                                                                               // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                                                 // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                                           // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                                                 // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                                                         // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [108:0] rsp_xbar_demux_002_src1_data;                                                                                                  // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	wire   [18:0] rsp_xbar_demux_002_src1_channel;                                                                                               // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                                                           // rsp_xbar_demux_003:src2_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                                                 // rsp_xbar_demux_003:src2_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                                                         // rsp_xbar_demux_003:src2_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire   [90:0] rsp_xbar_demux_003_src2_data;                                                                                                  // rsp_xbar_demux_003:src2_data -> rsp_xbar_mux_002:sink1_data
	wire   [18:0] rsp_xbar_demux_003_src2_channel;                                                                                               // rsp_xbar_demux_003:src2_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_003_src2_ready;                                                                                                 // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_003:src2_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                                           // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                                                 // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                                         // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	wire  [108:0] rsp_xbar_demux_004_src0_data;                                                                                                  // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src0_channel;                                                                                               // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                                                 // rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                                           // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                                                 // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                                         // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [108:0] rsp_xbar_demux_004_src1_data;                                                                                                  // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	wire   [18:0] rsp_xbar_demux_004_src1_channel;                                                                                               // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                                           // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux:sink5_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                                                 // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux:sink5_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                                         // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux:sink5_startofpacket
	wire  [108:0] rsp_xbar_demux_005_src0_data;                                                                                                  // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src0_channel;                                                                                               // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux:sink5_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                                                 // rsp_xbar_mux:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                                           // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                                                 // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_001:sink5_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                                         // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [108:0] rsp_xbar_demux_005_src1_data;                                                                                                  // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_001:sink5_data
	wire   [18:0] rsp_xbar_demux_005_src1_channel;                                                                                               // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_001:sink5_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                                           // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux:sink7_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                                                 // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux:sink7_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                                         // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux:sink7_startofpacket
	wire  [108:0] rsp_xbar_demux_007_src0_data;                                                                                                  // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src0_channel;                                                                                               // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux:sink7_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                                                 // rsp_xbar_mux:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_007_src1_endofpacket;                                                                                           // rsp_xbar_demux_007:src1_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          rsp_xbar_demux_007_src1_valid;                                                                                                 // rsp_xbar_demux_007:src1_valid -> rsp_xbar_mux_001:sink7_valid
	wire          rsp_xbar_demux_007_src1_startofpacket;                                                                                         // rsp_xbar_demux_007:src1_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [108:0] rsp_xbar_demux_007_src1_data;                                                                                                  // rsp_xbar_demux_007:src1_data -> rsp_xbar_mux_001:sink7_data
	wire   [18:0] rsp_xbar_demux_007_src1_channel;                                                                                               // rsp_xbar_demux_007:src1_channel -> rsp_xbar_mux_001:sink7_channel
	wire          rsp_xbar_demux_007_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src1_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                                           // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux:sink8_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                                                 // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux:sink8_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                                         // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux:sink8_startofpacket
	wire  [108:0] rsp_xbar_demux_008_src0_data;                                                                                                  // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux:sink8_data
	wire   [18:0] rsp_xbar_demux_008_src0_channel;                                                                                               // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux:sink8_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                                                 // rsp_xbar_mux:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                                           // rsp_xbar_demux_008:src1_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                                                 // rsp_xbar_demux_008:src1_valid -> rsp_xbar_mux_001:sink8_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                                                         // rsp_xbar_demux_008:src1_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [108:0] rsp_xbar_demux_008_src1_data;                                                                                                  // rsp_xbar_demux_008:src1_data -> rsp_xbar_mux_001:sink8_data
	wire   [18:0] rsp_xbar_demux_008_src1_channel;                                                                                               // rsp_xbar_demux_008:src1_channel -> rsp_xbar_mux_001:sink8_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src1_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                                           // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux:sink9_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                                                 // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux:sink9_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                                         // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux:sink9_startofpacket
	wire  [108:0] rsp_xbar_demux_009_src0_data;                                                                                                  // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src0_channel;                                                                                               // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux:sink9_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                                                 // rsp_xbar_mux:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                                           // rsp_xbar_demux_009:src1_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                                                 // rsp_xbar_demux_009:src1_valid -> rsp_xbar_mux_001:sink9_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                                                         // rsp_xbar_demux_009:src1_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [108:0] rsp_xbar_demux_009_src1_data;                                                                                                  // rsp_xbar_demux_009:src1_data -> rsp_xbar_mux_001:sink9_data
	wire   [18:0] rsp_xbar_demux_009_src1_channel;                                                                                               // rsp_xbar_demux_009:src1_channel -> rsp_xbar_mux_001:sink9_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src1_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                                           // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux:sink10_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                                                 // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux:sink10_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                                         // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux:sink10_startofpacket
	wire  [108:0] rsp_xbar_demux_010_src0_data;                                                                                                  // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src0_channel;                                                                                               // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux:sink10_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                                                 // rsp_xbar_mux:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                                           // rsp_xbar_demux_010:src1_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                                                 // rsp_xbar_demux_010:src1_valid -> rsp_xbar_mux_001:sink10_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                                                         // rsp_xbar_demux_010:src1_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [108:0] rsp_xbar_demux_010_src1_data;                                                                                                  // rsp_xbar_demux_010:src1_data -> rsp_xbar_mux_001:sink10_data
	wire   [18:0] rsp_xbar_demux_010_src1_channel;                                                                                               // rsp_xbar_demux_010:src1_channel -> rsp_xbar_mux_001:sink10_channel
	wire          rsp_xbar_demux_010_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src1_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                                           // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux:sink11_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                                                 // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux:sink11_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                                         // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux:sink11_startofpacket
	wire  [108:0] rsp_xbar_demux_011_src0_data;                                                                                                  // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux:sink11_data
	wire   [18:0] rsp_xbar_demux_011_src0_channel;                                                                                               // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux:sink11_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                                                 // rsp_xbar_mux:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_011_src1_endofpacket;                                                                                           // rsp_xbar_demux_011:src1_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire          rsp_xbar_demux_011_src1_valid;                                                                                                 // rsp_xbar_demux_011:src1_valid -> rsp_xbar_mux_001:sink11_valid
	wire          rsp_xbar_demux_011_src1_startofpacket;                                                                                         // rsp_xbar_demux_011:src1_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [108:0] rsp_xbar_demux_011_src1_data;                                                                                                  // rsp_xbar_demux_011:src1_data -> rsp_xbar_mux_001:sink11_data
	wire   [18:0] rsp_xbar_demux_011_src1_channel;                                                                                               // rsp_xbar_demux_011:src1_channel -> rsp_xbar_mux_001:sink11_channel
	wire          rsp_xbar_demux_011_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src1_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                                           // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux:sink12_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                                                 // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux:sink12_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                                         // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux:sink12_startofpacket
	wire  [108:0] rsp_xbar_demux_012_src0_data;                                                                                                  // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux:sink12_data
	wire   [18:0] rsp_xbar_demux_012_src0_channel;                                                                                               // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux:sink12_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                                                 // rsp_xbar_mux:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire          rsp_xbar_demux_012_src1_endofpacket;                                                                                           // rsp_xbar_demux_012:src1_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire          rsp_xbar_demux_012_src1_valid;                                                                                                 // rsp_xbar_demux_012:src1_valid -> rsp_xbar_mux_001:sink12_valid
	wire          rsp_xbar_demux_012_src1_startofpacket;                                                                                         // rsp_xbar_demux_012:src1_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [108:0] rsp_xbar_demux_012_src1_data;                                                                                                  // rsp_xbar_demux_012:src1_data -> rsp_xbar_mux_001:sink12_data
	wire   [18:0] rsp_xbar_demux_012_src1_channel;                                                                                               // rsp_xbar_demux_012:src1_channel -> rsp_xbar_mux_001:sink12_channel
	wire          rsp_xbar_demux_012_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src1_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                                           // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux:sink13_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                                                 // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux:sink13_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                                         // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux:sink13_startofpacket
	wire  [108:0] rsp_xbar_demux_013_src0_data;                                                                                                  // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux:sink13_data
	wire   [18:0] rsp_xbar_demux_013_src0_channel;                                                                                               // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux:sink13_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                                                 // rsp_xbar_mux:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire          rsp_xbar_demux_013_src1_endofpacket;                                                                                           // rsp_xbar_demux_013:src1_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire          rsp_xbar_demux_013_src1_valid;                                                                                                 // rsp_xbar_demux_013:src1_valid -> rsp_xbar_mux_001:sink13_valid
	wire          rsp_xbar_demux_013_src1_startofpacket;                                                                                         // rsp_xbar_demux_013:src1_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [108:0] rsp_xbar_demux_013_src1_data;                                                                                                  // rsp_xbar_demux_013:src1_data -> rsp_xbar_mux_001:sink13_data
	wire   [18:0] rsp_xbar_demux_013_src1_channel;                                                                                               // rsp_xbar_demux_013:src1_channel -> rsp_xbar_mux_001:sink13_channel
	wire          rsp_xbar_demux_013_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src1_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                                           // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux:sink14_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                                                 // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux:sink14_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                                         // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux:sink14_startofpacket
	wire  [108:0] rsp_xbar_demux_014_src0_data;                                                                                                  // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux:sink14_data
	wire   [18:0] rsp_xbar_demux_014_src0_channel;                                                                                               // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux:sink14_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                                                 // rsp_xbar_mux:sink14_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_014_src1_endofpacket;                                                                                           // rsp_xbar_demux_014:src1_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	wire          rsp_xbar_demux_014_src1_valid;                                                                                                 // rsp_xbar_demux_014:src1_valid -> rsp_xbar_mux_001:sink14_valid
	wire          rsp_xbar_demux_014_src1_startofpacket;                                                                                         // rsp_xbar_demux_014:src1_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	wire  [108:0] rsp_xbar_demux_014_src1_data;                                                                                                  // rsp_xbar_demux_014:src1_data -> rsp_xbar_mux_001:sink14_data
	wire   [18:0] rsp_xbar_demux_014_src1_channel;                                                                                               // rsp_xbar_demux_014:src1_channel -> rsp_xbar_mux_001:sink14_channel
	wire          rsp_xbar_demux_014_src1_ready;                                                                                                 // rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src1_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                                           // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                                                 // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                                         // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	wire  [108:0] rsp_xbar_demux_016_src0_data;                                                                                                  // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	wire   [18:0] rsp_xbar_demux_016_src0_channel;                                                                                               // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                                                 // rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                                           // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                                                 // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                                         // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	wire  [108:0] rsp_xbar_demux_017_src0_data;                                                                                                  // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	wire   [18:0] rsp_xbar_demux_017_src0_channel;                                                                                               // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                                                 // rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                                           // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                                                 // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                                         // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	wire  [108:0] rsp_xbar_demux_018_src0_data;                                                                                                  // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	wire   [18:0] rsp_xbar_demux_018_src0_channel;                                                                                               // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                                                 // rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                                                   // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                                                 // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [108:0] limiter_cmd_src_data;                                                                                                          // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire   [18:0] limiter_cmd_src_channel;                                                                                                       // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                                                         // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                                                  // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                                                        // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                                                // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [108:0] rsp_xbar_mux_src_data;                                                                                                         // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_src_channel;                                                                                                      // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                                                        // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                                               // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                                             // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [108:0] limiter_001_cmd_src_data;                                                                                                      // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire   [18:0] limiter_001_cmd_src_channel;                                                                                                   // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                                                     // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                                              // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                                                    // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                                            // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [108:0] rsp_xbar_mux_001_src_data;                                                                                                     // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire   [18:0] rsp_xbar_mux_001_src_channel;                                                                                                  // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                                                    // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          addr_router_002_src_endofpacket;                                                                                               // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                                                     // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                                             // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire   [90:0] addr_router_002_src_data;                                                                                                      // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire   [18:0] addr_router_002_src_channel;                                                                                                   // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                                                     // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                                              // rsp_xbar_mux_002:src_endofpacket -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                                                    // rsp_xbar_mux_002:src_valid -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                                            // rsp_xbar_mux_002:src_startofpacket -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [90:0] rsp_xbar_mux_002_src_data;                                                                                                     // rsp_xbar_mux_002:src_data -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire   [18:0] rsp_xbar_mux_002_src_channel;                                                                                                  // rsp_xbar_mux_002:src_channel -> amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                                                    // amd_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_002:src_ready
	wire          cmd_xbar_mux_src_endofpacket;                                                                                                  // cmd_xbar_mux:src_endofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                                        // cmd_xbar_mux:src_valid -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                                                // cmd_xbar_mux:src_startofpacket -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_src_data;                                                                                                         // cmd_xbar_mux:src_data -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_src_channel;                                                                                                      // cmd_xbar_mux:src_channel -> nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                                        // nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                                                     // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                                           // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                                                   // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [108:0] id_router_src_data;                                                                                                            // id_router:src_data -> rsp_xbar_demux:sink_data
	wire   [18:0] id_router_src_channel;                                                                                                         // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                                           // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                                              // cmd_xbar_mux_001:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                                                    // cmd_xbar_mux_001:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                                            // cmd_xbar_mux_001:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_001_src_data;                                                                                                     // cmd_xbar_mux_001:src_data -> burst_adapter:sink0_data
	wire   [18:0] cmd_xbar_mux_001_src_channel;                                                                                                  // cmd_xbar_mux_001:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                                                    // burst_adapter:sink0_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                                                 // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                                       // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                                               // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire   [90:0] id_router_001_src_data;                                                                                                        // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire   [18:0] id_router_001_src_channel;                                                                                                     // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                                       // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                                              // cmd_xbar_mux_002:src_endofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                                                    // cmd_xbar_mux_002:src_valid -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                                            // cmd_xbar_mux_002:src_startofpacket -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_002_src_data;                                                                                                     // cmd_xbar_mux_002:src_data -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_002_src_channel;                                                                                                  // cmd_xbar_mux_002:src_channel -> onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                                                    // onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                                                 // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                                       // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                                               // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [108:0] id_router_002_src_data;                                                                                                        // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire   [18:0] id_router_002_src_channel;                                                                                                     // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                                       // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                                              // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                                                    // cmd_xbar_mux_003:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                                            // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_003_src_data;                                                                                                     // cmd_xbar_mux_003:src_data -> burst_adapter_001:sink0_data
	wire   [18:0] cmd_xbar_mux_003_src_channel;                                                                                                  // cmd_xbar_mux_003:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                                                    // burst_adapter_001:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                                                 // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                                       // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                                               // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire   [90:0] id_router_003_src_data;                                                                                                        // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire   [18:0] id_router_003_src_channel;                                                                                                     // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                                       // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                                              // cmd_xbar_mux_004:src_endofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                                                    // cmd_xbar_mux_004:src_valid -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                                            // cmd_xbar_mux_004:src_startofpacket -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_004_src_data;                                                                                                     // cmd_xbar_mux_004:src_data -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_004_src_channel;                                                                                                  // cmd_xbar_mux_004:src_channel -> rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                                                    // rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                                                 // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                                       // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                                               // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [108:0] id_router_004_src_data;                                                                                                        // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire   [18:0] id_router_004_src_channel;                                                                                                     // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                                       // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                                              // cmd_xbar_mux_005:src_endofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                                                    // cmd_xbar_mux_005:src_valid -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                                            // cmd_xbar_mux_005:src_startofpacket -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_005_src_data;                                                                                                     // cmd_xbar_mux_005:src_data -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_005_src_channel;                                                                                                  // cmd_xbar_mux_005:src_channel -> pio_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                                                    // pio_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                                                 // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                                       // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                                               // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [108:0] id_router_005_src_data;                                                                                                        // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire   [18:0] id_router_005_src_channel;                                                                                                     // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                                       // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                                              // cmd_xbar_mux_006:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                                                    // cmd_xbar_mux_006:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                                                            // cmd_xbar_mux_006:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire   [81:0] cmd_xbar_mux_006_src_data;                                                                                                     // cmd_xbar_mux_006:src_data -> burst_adapter_002:sink0_data
	wire   [18:0] cmd_xbar_mux_006_src_channel;                                                                                                  // cmd_xbar_mux_006:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                                                    // burst_adapter_002:sink0_ready -> cmd_xbar_mux_006:src_ready
	wire          id_router_006_src_endofpacket;                                                                                                 // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                                       // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                                               // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire   [81:0] id_router_006_src_data;                                                                                                        // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire   [18:0] id_router_006_src_channel;                                                                                                     // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                                       // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_mux_007_src_endofpacket;                                                                                              // cmd_xbar_mux_007:src_endofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_007_src_valid;                                                                                                    // cmd_xbar_mux_007:src_valid -> pio_3_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_007_src_startofpacket;                                                                                            // cmd_xbar_mux_007:src_startofpacket -> pio_3_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_007_src_data;                                                                                                     // cmd_xbar_mux_007:src_data -> pio_3_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_007_src_channel;                                                                                                  // cmd_xbar_mux_007:src_channel -> pio_3_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_007_src_ready;                                                                                                    // pio_3_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_007:src_ready
	wire          id_router_007_src_endofpacket;                                                                                                 // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                                       // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                                               // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [108:0] id_router_007_src_data;                                                                                                        // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [18:0] id_router_007_src_channel;                                                                                                     // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                                       // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                                              // cmd_xbar_mux_008:src_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                                                    // cmd_xbar_mux_008:src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                                            // cmd_xbar_mux_008:src_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_008_src_data;                                                                                                     // cmd_xbar_mux_008:src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_008_src_channel;                                                                                                  // cmd_xbar_mux_008:src_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                                                 // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                                       // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                                               // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [108:0] id_router_008_src_data;                                                                                                        // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [18:0] id_router_008_src_channel;                                                                                                     // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                                       // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                                              // cmd_xbar_mux_009:src_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                                                    // cmd_xbar_mux_009:src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                                            // cmd_xbar_mux_009:src_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_009_src_data;                                                                                                     // cmd_xbar_mux_009:src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_009_src_channel;                                                                                                  // cmd_xbar_mux_009:src_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                                                    // timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                                                 // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                                       // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                                               // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [108:0] id_router_009_src_data;                                                                                                        // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [18:0] id_router_009_src_channel;                                                                                                     // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                                       // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                                              // cmd_xbar_mux_010:src_endofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                                                    // cmd_xbar_mux_010:src_valid -> pio_4_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                                            // cmd_xbar_mux_010:src_startofpacket -> pio_4_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_010_src_data;                                                                                                     // cmd_xbar_mux_010:src_data -> pio_4_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_010_src_channel;                                                                                                  // cmd_xbar_mux_010:src_channel -> pio_4_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                                                    // pio_4_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_010:src_ready
	wire          id_router_010_src_endofpacket;                                                                                                 // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                                       // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                                               // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [108:0] id_router_010_src_data;                                                                                                        // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [18:0] id_router_010_src_channel;                                                                                                     // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                                       // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_mux_011_src_endofpacket;                                                                                              // cmd_xbar_mux_011:src_endofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_011_src_valid;                                                                                                    // cmd_xbar_mux_011:src_valid -> pio_5_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_011_src_startofpacket;                                                                                            // cmd_xbar_mux_011:src_startofpacket -> pio_5_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_011_src_data;                                                                                                     // cmd_xbar_mux_011:src_data -> pio_5_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_011_src_channel;                                                                                                  // cmd_xbar_mux_011:src_channel -> pio_5_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_011_src_ready;                                                                                                    // pio_5_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_011:src_ready
	wire          id_router_011_src_endofpacket;                                                                                                 // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                                       // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                                               // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [108:0] id_router_011_src_data;                                                                                                        // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [18:0] id_router_011_src_channel;                                                                                                     // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                                       // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          cmd_xbar_mux_012_src_endofpacket;                                                                                              // cmd_xbar_mux_012:src_endofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_012_src_valid;                                                                                                    // cmd_xbar_mux_012:src_valid -> pio_6_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_012_src_startofpacket;                                                                                            // cmd_xbar_mux_012:src_startofpacket -> pio_6_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_012_src_data;                                                                                                     // cmd_xbar_mux_012:src_data -> pio_6_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_012_src_channel;                                                                                                  // cmd_xbar_mux_012:src_channel -> pio_6_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_012_src_ready;                                                                                                    // pio_6_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_012:src_ready
	wire          id_router_012_src_endofpacket;                                                                                                 // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                                       // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                                               // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [108:0] id_router_012_src_data;                                                                                                        // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [18:0] id_router_012_src_channel;                                                                                                     // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                                       // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          cmd_xbar_mux_013_src_endofpacket;                                                                                              // cmd_xbar_mux_013:src_endofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_013_src_valid;                                                                                                    // cmd_xbar_mux_013:src_valid -> pio_7_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_013_src_startofpacket;                                                                                            // cmd_xbar_mux_013:src_startofpacket -> pio_7_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_013_src_data;                                                                                                     // cmd_xbar_mux_013:src_data -> pio_7_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_013_src_channel;                                                                                                  // cmd_xbar_mux_013:src_channel -> pio_7_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_013_src_ready;                                                                                                    // pio_7_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_013:src_ready
	wire          id_router_013_src_endofpacket;                                                                                                 // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                                       // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                                               // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [108:0] id_router_013_src_data;                                                                                                        // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [18:0] id_router_013_src_channel;                                                                                                     // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                                       // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_mux_014_src_endofpacket;                                                                                              // cmd_xbar_mux_014:src_endofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_014_src_valid;                                                                                                    // cmd_xbar_mux_014:src_valid -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_014_src_startofpacket;                                                                                            // cmd_xbar_mux_014:src_startofpacket -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [108:0] cmd_xbar_mux_014_src_data;                                                                                                     // cmd_xbar_mux_014:src_data -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [18:0] cmd_xbar_mux_014_src_channel;                                                                                                  // cmd_xbar_mux_014:src_channel -> Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_014_src_ready;                                                                                                    // Altera_UP_SD_Card_Avalon_Interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_014:src_ready
	wire          id_router_014_src_endofpacket;                                                                                                 // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                                       // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                                               // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire  [108:0] id_router_014_src_data;                                                                                                        // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [18:0] id_router_014_src_channel;                                                                                                     // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                                       // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_mux_015_src_endofpacket;                                                                                              // cmd_xbar_mux_015:src_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_mux_015_src_valid;                                                                                                    // cmd_xbar_mux_015:src_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_mux_015_src_startofpacket;                                                                                            // cmd_xbar_mux_015:src_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire   [90:0] cmd_xbar_mux_015_src_data;                                                                                                     // cmd_xbar_mux_015:src_data -> burst_adapter_003:sink0_data
	wire   [18:0] cmd_xbar_mux_015_src_channel;                                                                                                  // cmd_xbar_mux_015:src_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_mux_015_src_ready;                                                                                                    // burst_adapter_003:sink0_ready -> cmd_xbar_mux_015:src_ready
	wire          id_router_015_src_endofpacket;                                                                                                 // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                                       // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                                               // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [90:0] id_router_015_src_data;                                                                                                        // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [18:0] id_router_015_src_channel;                                                                                                     // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                                       // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_001_src16_ready;                                                                                                // jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	wire          id_router_016_src_endofpacket;                                                                                                 // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                                       // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                                               // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire  [108:0] id_router_016_src_data;                                                                                                        // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [18:0] id_router_016_src_channel;                                                                                                     // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                                       // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_001_src17_ready;                                                                                                // pio_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	wire          id_router_017_src_endofpacket;                                                                                                 // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                                       // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                                               // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire  [108:0] id_router_017_src_data;                                                                                                        // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [18:0] id_router_017_src_channel;                                                                                                     // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                                       // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_001_src18_ready;                                                                                                // pio_2_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	wire          id_router_018_src_endofpacket;                                                                                                 // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                                       // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                                               // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire  [108:0] id_router_018_src_data;                                                                                                        // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire   [18:0] id_router_018_src_channel;                                                                                                     // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                                       // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_src1_endofpacket;                                                                                               // cmd_xbar_demux:src1_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                                                     // cmd_xbar_demux:src1_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                                             // cmd_xbar_demux:src1_startofpacket -> width_adapter:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src1_data;                                                                                                      // cmd_xbar_demux:src1_data -> width_adapter:in_data
	wire   [18:0] cmd_xbar_demux_src1_channel;                                                                                                   // cmd_xbar_demux:src1_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_ready;                                                                                                     // width_adapter:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_src_endofpacket;                                                                                                 // width_adapter:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                                                       // width_adapter:out_valid -> cmd_xbar_mux_001:sink0_valid
	wire          width_adapter_src_startofpacket;                                                                                               // width_adapter:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire   [90:0] width_adapter_src_data;                                                                                                        // width_adapter:out_data -> cmd_xbar_mux_001:sink0_data
	wire          width_adapter_src_ready;                                                                                                       // cmd_xbar_mux_001:sink0_ready -> width_adapter:out_ready
	wire   [18:0] width_adapter_src_channel;                                                                                                     // width_adapter:out_channel -> cmd_xbar_mux_001:sink0_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                                                               // cmd_xbar_demux:src3_endofpacket -> width_adapter_001:in_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                                                                     // cmd_xbar_demux:src3_valid -> width_adapter_001:in_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                                                             // cmd_xbar_demux:src3_startofpacket -> width_adapter_001:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src3_data;                                                                                                      // cmd_xbar_demux:src3_data -> width_adapter_001:in_data
	wire   [18:0] cmd_xbar_demux_src3_channel;                                                                                                   // cmd_xbar_demux:src3_channel -> width_adapter_001:in_channel
	wire          cmd_xbar_demux_src3_ready;                                                                                                     // width_adapter_001:in_ready -> cmd_xbar_demux:src3_ready
	wire          width_adapter_001_src_endofpacket;                                                                                             // width_adapter_001:out_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          width_adapter_001_src_valid;                                                                                                   // width_adapter_001:out_valid -> cmd_xbar_mux_003:sink0_valid
	wire          width_adapter_001_src_startofpacket;                                                                                           // width_adapter_001:out_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire   [90:0] width_adapter_001_src_data;                                                                                                    // width_adapter_001:out_data -> cmd_xbar_mux_003:sink0_data
	wire          width_adapter_001_src_ready;                                                                                                   // cmd_xbar_mux_003:sink0_ready -> width_adapter_001:out_ready
	wire   [18:0] width_adapter_001_src_channel;                                                                                                 // width_adapter_001:out_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_src6_endofpacket;                                                                                               // cmd_xbar_demux:src6_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_src6_valid;                                                                                                     // cmd_xbar_demux:src6_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_src6_startofpacket;                                                                                             // cmd_xbar_demux:src6_startofpacket -> width_adapter_002:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src6_data;                                                                                                      // cmd_xbar_demux:src6_data -> width_adapter_002:in_data
	wire   [18:0] cmd_xbar_demux_src6_channel;                                                                                                   // cmd_xbar_demux:src6_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_src6_ready;                                                                                                     // width_adapter_002:in_ready -> cmd_xbar_demux:src6_ready
	wire          width_adapter_002_src_endofpacket;                                                                                             // width_adapter_002:out_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                                                                   // width_adapter_002:out_valid -> cmd_xbar_mux_006:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                                                           // width_adapter_002:out_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire   [81:0] width_adapter_002_src_data;                                                                                                    // width_adapter_002:out_data -> cmd_xbar_mux_006:sink0_data
	wire          width_adapter_002_src_ready;                                                                                                   // cmd_xbar_mux_006:sink0_ready -> width_adapter_002:out_ready
	wire   [18:0] width_adapter_002_src_channel;                                                                                                 // width_adapter_002:out_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_src15_endofpacket;                                                                                              // cmd_xbar_demux:src15_endofpacket -> width_adapter_003:in_endofpacket
	wire          cmd_xbar_demux_src15_valid;                                                                                                    // cmd_xbar_demux:src15_valid -> width_adapter_003:in_valid
	wire          cmd_xbar_demux_src15_startofpacket;                                                                                            // cmd_xbar_demux:src15_startofpacket -> width_adapter_003:in_startofpacket
	wire  [108:0] cmd_xbar_demux_src15_data;                                                                                                     // cmd_xbar_demux:src15_data -> width_adapter_003:in_data
	wire   [18:0] cmd_xbar_demux_src15_channel;                                                                                                  // cmd_xbar_demux:src15_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_demux_src15_ready;                                                                                                    // width_adapter_003:in_ready -> cmd_xbar_demux:src15_ready
	wire          width_adapter_003_src_endofpacket;                                                                                             // width_adapter_003:out_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	wire          width_adapter_003_src_valid;                                                                                                   // width_adapter_003:out_valid -> cmd_xbar_mux_015:sink0_valid
	wire          width_adapter_003_src_startofpacket;                                                                                           // width_adapter_003:out_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	wire   [90:0] width_adapter_003_src_data;                                                                                                    // width_adapter_003:out_data -> cmd_xbar_mux_015:sink0_data
	wire          width_adapter_003_src_ready;                                                                                                   // cmd_xbar_mux_015:sink0_ready -> width_adapter_003:out_ready
	wire   [18:0] width_adapter_003_src_channel;                                                                                                 // width_adapter_003:out_channel -> cmd_xbar_mux_015:sink0_channel
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                                           // cmd_xbar_demux_001:src1_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                                                 // cmd_xbar_demux_001:src1_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                                                         // cmd_xbar_demux_001:src1_startofpacket -> width_adapter_004:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src1_data;                                                                                                  // cmd_xbar_demux_001:src1_data -> width_adapter_004:in_data
	wire   [18:0] cmd_xbar_demux_001_src1_channel;                                                                                               // cmd_xbar_demux_001:src1_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                                                 // width_adapter_004:in_ready -> cmd_xbar_demux_001:src1_ready
	wire          width_adapter_004_src_endofpacket;                                                                                             // width_adapter_004:out_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_004_src_valid;                                                                                                   // width_adapter_004:out_valid -> cmd_xbar_mux_001:sink1_valid
	wire          width_adapter_004_src_startofpacket;                                                                                           // width_adapter_004:out_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire   [90:0] width_adapter_004_src_data;                                                                                                    // width_adapter_004:out_data -> cmd_xbar_mux_001:sink1_data
	wire          width_adapter_004_src_ready;                                                                                                   // cmd_xbar_mux_001:sink1_ready -> width_adapter_004:out_ready
	wire   [18:0] width_adapter_004_src_channel;                                                                                                 // width_adapter_004:out_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                                           // cmd_xbar_demux_001:src3_endofpacket -> width_adapter_005:in_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                                                 // cmd_xbar_demux_001:src3_valid -> width_adapter_005:in_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                                                         // cmd_xbar_demux_001:src3_startofpacket -> width_adapter_005:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src3_data;                                                                                                  // cmd_xbar_demux_001:src3_data -> width_adapter_005:in_data
	wire   [18:0] cmd_xbar_demux_001_src3_channel;                                                                                               // cmd_xbar_demux_001:src3_channel -> width_adapter_005:in_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                                                 // width_adapter_005:in_ready -> cmd_xbar_demux_001:src3_ready
	wire          width_adapter_005_src_endofpacket;                                                                                             // width_adapter_005:out_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          width_adapter_005_src_valid;                                                                                                   // width_adapter_005:out_valid -> cmd_xbar_mux_003:sink1_valid
	wire          width_adapter_005_src_startofpacket;                                                                                           // width_adapter_005:out_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire   [90:0] width_adapter_005_src_data;                                                                                                    // width_adapter_005:out_data -> cmd_xbar_mux_003:sink1_data
	wire          width_adapter_005_src_ready;                                                                                                   // cmd_xbar_mux_003:sink1_ready -> width_adapter_005:out_ready
	wire   [18:0] width_adapter_005_src_channel;                                                                                                 // width_adapter_005:out_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                                           // cmd_xbar_demux_001:src6_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                                                 // cmd_xbar_demux_001:src6_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                                                         // cmd_xbar_demux_001:src6_startofpacket -> width_adapter_006:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src6_data;                                                                                                  // cmd_xbar_demux_001:src6_data -> width_adapter_006:in_data
	wire   [18:0] cmd_xbar_demux_001_src6_channel;                                                                                               // cmd_xbar_demux_001:src6_channel -> width_adapter_006:in_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                                                 // width_adapter_006:in_ready -> cmd_xbar_demux_001:src6_ready
	wire          width_adapter_006_src_endofpacket;                                                                                             // width_adapter_006:out_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          width_adapter_006_src_valid;                                                                                                   // width_adapter_006:out_valid -> cmd_xbar_mux_006:sink1_valid
	wire          width_adapter_006_src_startofpacket;                                                                                           // width_adapter_006:out_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire   [81:0] width_adapter_006_src_data;                                                                                                    // width_adapter_006:out_data -> cmd_xbar_mux_006:sink1_data
	wire          width_adapter_006_src_ready;                                                                                                   // cmd_xbar_mux_006:sink1_ready -> width_adapter_006:out_ready
	wire   [18:0] width_adapter_006_src_channel;                                                                                                 // width_adapter_006:out_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_001_src15_endofpacket;                                                                                          // cmd_xbar_demux_001:src15_endofpacket -> width_adapter_007:in_endofpacket
	wire          cmd_xbar_demux_001_src15_valid;                                                                                                // cmd_xbar_demux_001:src15_valid -> width_adapter_007:in_valid
	wire          cmd_xbar_demux_001_src15_startofpacket;                                                                                        // cmd_xbar_demux_001:src15_startofpacket -> width_adapter_007:in_startofpacket
	wire  [108:0] cmd_xbar_demux_001_src15_data;                                                                                                 // cmd_xbar_demux_001:src15_data -> width_adapter_007:in_data
	wire   [18:0] cmd_xbar_demux_001_src15_channel;                                                                                              // cmd_xbar_demux_001:src15_channel -> width_adapter_007:in_channel
	wire          cmd_xbar_demux_001_src15_ready;                                                                                                // width_adapter_007:in_ready -> cmd_xbar_demux_001:src15_ready
	wire          width_adapter_007_src_endofpacket;                                                                                             // width_adapter_007:out_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	wire          width_adapter_007_src_valid;                                                                                                   // width_adapter_007:out_valid -> cmd_xbar_mux_015:sink1_valid
	wire          width_adapter_007_src_startofpacket;                                                                                           // width_adapter_007:out_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	wire   [90:0] width_adapter_007_src_data;                                                                                                    // width_adapter_007:out_data -> cmd_xbar_mux_015:sink1_data
	wire          width_adapter_007_src_ready;                                                                                                   // cmd_xbar_mux_015:sink1_ready -> width_adapter_007:out_ready
	wire   [18:0] width_adapter_007_src_channel;                                                                                                 // width_adapter_007:out_channel -> cmd_xbar_mux_015:sink1_channel
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                                           // rsp_xbar_demux_001:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                                                 // rsp_xbar_demux_001:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                                         // rsp_xbar_demux_001:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src0_data;                                                                                                  // rsp_xbar_demux_001:src0_data -> width_adapter_008:in_data
	wire   [18:0] rsp_xbar_demux_001_src0_channel;                                                                                               // rsp_xbar_demux_001:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                                                 // width_adapter_008:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                                             // width_adapter_008:out_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          width_adapter_008_src_valid;                                                                                                   // width_adapter_008:out_valid -> rsp_xbar_mux:sink1_valid
	wire          width_adapter_008_src_startofpacket;                                                                                           // width_adapter_008:out_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [108:0] width_adapter_008_src_data;                                                                                                    // width_adapter_008:out_data -> rsp_xbar_mux:sink1_data
	wire          width_adapter_008_src_ready;                                                                                                   // rsp_xbar_mux:sink1_ready -> width_adapter_008:out_ready
	wire   [18:0] width_adapter_008_src_channel;                                                                                                 // width_adapter_008:out_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                                           // rsp_xbar_demux_001:src1_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                                                 // rsp_xbar_demux_001:src1_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                                         // rsp_xbar_demux_001:src1_startofpacket -> width_adapter_009:in_startofpacket
	wire   [90:0] rsp_xbar_demux_001_src1_data;                                                                                                  // rsp_xbar_demux_001:src1_data -> width_adapter_009:in_data
	wire   [18:0] rsp_xbar_demux_001_src1_channel;                                                                                               // rsp_xbar_demux_001:src1_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                                                 // width_adapter_009:in_ready -> rsp_xbar_demux_001:src1_ready
	wire          width_adapter_009_src_endofpacket;                                                                                             // width_adapter_009:out_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          width_adapter_009_src_valid;                                                                                                   // width_adapter_009:out_valid -> rsp_xbar_mux_001:sink1_valid
	wire          width_adapter_009_src_startofpacket;                                                                                           // width_adapter_009:out_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [108:0] width_adapter_009_src_data;                                                                                                    // width_adapter_009:out_data -> rsp_xbar_mux_001:sink1_data
	wire          width_adapter_009_src_ready;                                                                                                   // rsp_xbar_mux_001:sink1_ready -> width_adapter_009:out_ready
	wire   [18:0] width_adapter_009_src_channel;                                                                                                 // width_adapter_009:out_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                                           // rsp_xbar_demux_003:src0_endofpacket -> width_adapter_010:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                                                 // rsp_xbar_demux_003:src0_valid -> width_adapter_010:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                                         // rsp_xbar_demux_003:src0_startofpacket -> width_adapter_010:in_startofpacket
	wire   [90:0] rsp_xbar_demux_003_src0_data;                                                                                                  // rsp_xbar_demux_003:src0_data -> width_adapter_010:in_data
	wire   [18:0] rsp_xbar_demux_003_src0_channel;                                                                                               // rsp_xbar_demux_003:src0_channel -> width_adapter_010:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                                                 // width_adapter_010:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          width_adapter_010_src_endofpacket;                                                                                             // width_adapter_010:out_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          width_adapter_010_src_valid;                                                                                                   // width_adapter_010:out_valid -> rsp_xbar_mux:sink3_valid
	wire          width_adapter_010_src_startofpacket;                                                                                           // width_adapter_010:out_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [108:0] width_adapter_010_src_data;                                                                                                    // width_adapter_010:out_data -> rsp_xbar_mux:sink3_data
	wire          width_adapter_010_src_ready;                                                                                                   // rsp_xbar_mux:sink3_ready -> width_adapter_010:out_ready
	wire   [18:0] width_adapter_010_src_channel;                                                                                                 // width_adapter_010:out_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                                           // rsp_xbar_demux_003:src1_endofpacket -> width_adapter_011:in_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                                                 // rsp_xbar_demux_003:src1_valid -> width_adapter_011:in_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                                         // rsp_xbar_demux_003:src1_startofpacket -> width_adapter_011:in_startofpacket
	wire   [90:0] rsp_xbar_demux_003_src1_data;                                                                                                  // rsp_xbar_demux_003:src1_data -> width_adapter_011:in_data
	wire   [18:0] rsp_xbar_demux_003_src1_channel;                                                                                               // rsp_xbar_demux_003:src1_channel -> width_adapter_011:in_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                                                 // width_adapter_011:in_ready -> rsp_xbar_demux_003:src1_ready
	wire          width_adapter_011_src_endofpacket;                                                                                             // width_adapter_011:out_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          width_adapter_011_src_valid;                                                                                                   // width_adapter_011:out_valid -> rsp_xbar_mux_001:sink3_valid
	wire          width_adapter_011_src_startofpacket;                                                                                           // width_adapter_011:out_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [108:0] width_adapter_011_src_data;                                                                                                    // width_adapter_011:out_data -> rsp_xbar_mux_001:sink3_data
	wire          width_adapter_011_src_ready;                                                                                                   // rsp_xbar_mux_001:sink3_ready -> width_adapter_011:out_ready
	wire   [18:0] width_adapter_011_src_channel;                                                                                                 // width_adapter_011:out_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                                           // rsp_xbar_demux_006:src0_endofpacket -> width_adapter_012:in_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                                                 // rsp_xbar_demux_006:src0_valid -> width_adapter_012:in_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                                         // rsp_xbar_demux_006:src0_startofpacket -> width_adapter_012:in_startofpacket
	wire   [81:0] rsp_xbar_demux_006_src0_data;                                                                                                  // rsp_xbar_demux_006:src0_data -> width_adapter_012:in_data
	wire   [18:0] rsp_xbar_demux_006_src0_channel;                                                                                               // rsp_xbar_demux_006:src0_channel -> width_adapter_012:in_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                                                 // width_adapter_012:in_ready -> rsp_xbar_demux_006:src0_ready
	wire          width_adapter_012_src_endofpacket;                                                                                             // width_adapter_012:out_endofpacket -> rsp_xbar_mux:sink6_endofpacket
	wire          width_adapter_012_src_valid;                                                                                                   // width_adapter_012:out_valid -> rsp_xbar_mux:sink6_valid
	wire          width_adapter_012_src_startofpacket;                                                                                           // width_adapter_012:out_startofpacket -> rsp_xbar_mux:sink6_startofpacket
	wire  [108:0] width_adapter_012_src_data;                                                                                                    // width_adapter_012:out_data -> rsp_xbar_mux:sink6_data
	wire          width_adapter_012_src_ready;                                                                                                   // rsp_xbar_mux:sink6_ready -> width_adapter_012:out_ready
	wire   [18:0] width_adapter_012_src_channel;                                                                                                 // width_adapter_012:out_channel -> rsp_xbar_mux:sink6_channel
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                                                           // rsp_xbar_demux_006:src1_endofpacket -> width_adapter_013:in_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                                                 // rsp_xbar_demux_006:src1_valid -> width_adapter_013:in_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                                                         // rsp_xbar_demux_006:src1_startofpacket -> width_adapter_013:in_startofpacket
	wire   [81:0] rsp_xbar_demux_006_src1_data;                                                                                                  // rsp_xbar_demux_006:src1_data -> width_adapter_013:in_data
	wire   [18:0] rsp_xbar_demux_006_src1_channel;                                                                                               // rsp_xbar_demux_006:src1_channel -> width_adapter_013:in_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                                                 // width_adapter_013:in_ready -> rsp_xbar_demux_006:src1_ready
	wire          width_adapter_013_src_endofpacket;                                                                                             // width_adapter_013:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          width_adapter_013_src_valid;                                                                                                   // width_adapter_013:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire          width_adapter_013_src_startofpacket;                                                                                           // width_adapter_013:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [108:0] width_adapter_013_src_data;                                                                                                    // width_adapter_013:out_data -> rsp_xbar_mux_001:sink6_data
	wire          width_adapter_013_src_ready;                                                                                                   // rsp_xbar_mux_001:sink6_ready -> width_adapter_013:out_ready
	wire   [18:0] width_adapter_013_src_channel;                                                                                                 // width_adapter_013:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                                           // rsp_xbar_demux_015:src0_endofpacket -> width_adapter_014:in_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                                                 // rsp_xbar_demux_015:src0_valid -> width_adapter_014:in_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                                         // rsp_xbar_demux_015:src0_startofpacket -> width_adapter_014:in_startofpacket
	wire   [90:0] rsp_xbar_demux_015_src0_data;                                                                                                  // rsp_xbar_demux_015:src0_data -> width_adapter_014:in_data
	wire   [18:0] rsp_xbar_demux_015_src0_channel;                                                                                               // rsp_xbar_demux_015:src0_channel -> width_adapter_014:in_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                                                 // width_adapter_014:in_ready -> rsp_xbar_demux_015:src0_ready
	wire          width_adapter_014_src_endofpacket;                                                                                             // width_adapter_014:out_endofpacket -> rsp_xbar_mux:sink15_endofpacket
	wire          width_adapter_014_src_valid;                                                                                                   // width_adapter_014:out_valid -> rsp_xbar_mux:sink15_valid
	wire          width_adapter_014_src_startofpacket;                                                                                           // width_adapter_014:out_startofpacket -> rsp_xbar_mux:sink15_startofpacket
	wire  [108:0] width_adapter_014_src_data;                                                                                                    // width_adapter_014:out_data -> rsp_xbar_mux:sink15_data
	wire          width_adapter_014_src_ready;                                                                                                   // rsp_xbar_mux:sink15_ready -> width_adapter_014:out_ready
	wire   [18:0] width_adapter_014_src_channel;                                                                                                 // width_adapter_014:out_channel -> rsp_xbar_mux:sink15_channel
	wire          rsp_xbar_demux_015_src1_endofpacket;                                                                                           // rsp_xbar_demux_015:src1_endofpacket -> width_adapter_015:in_endofpacket
	wire          rsp_xbar_demux_015_src1_valid;                                                                                                 // rsp_xbar_demux_015:src1_valid -> width_adapter_015:in_valid
	wire          rsp_xbar_demux_015_src1_startofpacket;                                                                                         // rsp_xbar_demux_015:src1_startofpacket -> width_adapter_015:in_startofpacket
	wire   [90:0] rsp_xbar_demux_015_src1_data;                                                                                                  // rsp_xbar_demux_015:src1_data -> width_adapter_015:in_data
	wire   [18:0] rsp_xbar_demux_015_src1_channel;                                                                                               // rsp_xbar_demux_015:src1_channel -> width_adapter_015:in_channel
	wire          rsp_xbar_demux_015_src1_ready;                                                                                                 // width_adapter_015:in_ready -> rsp_xbar_demux_015:src1_ready
	wire          width_adapter_015_src_endofpacket;                                                                                             // width_adapter_015:out_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	wire          width_adapter_015_src_valid;                                                                                                   // width_adapter_015:out_valid -> rsp_xbar_mux_001:sink15_valid
	wire          width_adapter_015_src_startofpacket;                                                                                           // width_adapter_015:out_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	wire  [108:0] width_adapter_015_src_data;                                                                                                    // width_adapter_015:out_data -> rsp_xbar_mux_001:sink15_data
	wire          width_adapter_015_src_ready;                                                                                                   // rsp_xbar_mux_001:sink15_ready -> width_adapter_015:out_ready
	wire   [18:0] width_adapter_015_src_channel;                                                                                                 // width_adapter_015:out_channel -> rsp_xbar_mux_001:sink15_channel
	wire   [18:0] limiter_cmd_valid_data;                                                                                                        // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [18:0] limiter_001_cmd_valid_data;                                                                                                    // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                                                      // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                                                      // to_external_bus_bridge_0:avalon_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                                                      // rs232_0:irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                                                                      // timer_0:irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                                                                                      // timer_1:irq -> irq_mapper:receiver4_irq
	wire   [31:0] nios2_qsys_0_d_irq_irq;                                                                                                        // irq_mapper:sender_irq -> nios2_qsys_0:d_irq

	nios_system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (up_clocks_0_sys_clk_clk),                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_0_data_master_address),                                          //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                             //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                                            //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                                      //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	nios_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (up_clocks_0_sys_clk_clk),                                       //   clk1.clk
		.address    (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.clken      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.chipselect (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.write      (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),      //       .write
		.readdata   (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.writedata  (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                             //       .reset_req
	);

	nios_system_jtag_uart_0 jtag_uart_0 (
		.clk            (up_clocks_0_sys_clk_clk),                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                          //             reset.reset_n
		.av_chipselect  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                  //               irq.irq
	);

	nios_system_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (up_clocks_0_sys_clk_clk),                                                //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                                        // reset.reset_n
		.az_addr        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                                        //  wire.export
		.zs_ba          (sdram_wire_ba),                                                          //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                                       //      .export
		.zs_cke         (sdram_wire_cke),                                                         //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                                        //      .export
		.zs_dq          (sdram_wire_dq),                                                          //      .export
		.zs_dqm         (sdram_wire_dqm),                                                         //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                                       //      .export
		.zs_we_n        (sdram_wire_we_n)                                                         //      .export
	);

	nios_system_up_clocks_0 up_clocks_0 (
		.CLOCK_50    (clk_clk),                            //       clk_in_primary.clk
		.reset       (rst_controller_001_reset_out_reset), // clk_in_primary_reset.reset
		.sys_clk     (up_clocks_0_sys_clk_clk),            //              sys_clk.clk
		.sys_reset_n (),                                   //        sys_clk_reset.reset_n
		.SDRAM_CLK   (sdram_clk_clk)                       //            sdram_clk.clk
	);

	nios_system_to_external_bus_bridge_0 to_external_bus_bridge_0 (
		.clk                (up_clocks_0_sys_clk_clk),                                                          //        clock_reset.clk
		.reset              (rst_controller_reset_out_reset),                                                   //  clock_reset_reset.reset
		.avalon_address     (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_address),     //       avalon_slave.address
		.avalon_byteenable  (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_byteenable),  //                   .byteenable
		.avalon_chipselect  (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.avalon_read        (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.avalon_write       (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.avalon_writedata   (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.avalon_readdata    (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.avalon_waitrequest (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.avalon_irq         (irq_mapper_receiver1_irq),                                                         //          interrupt.irq
		.acknowledge        (io_acknowledge),                                                                   // external_interface.export
		.irq                (io_irq),                                                                           //                   .export
		.address            (io_address),                                                                       //                   .export
		.bus_enable         (io_bus_enable),                                                                    //                   .export
		.byte_enable        (io_byte_enable),                                                                   //                   .export
		.rw                 (io_rw),                                                                            //                   .export
		.write_data         (io_write_data),                                                                    //                   .export
		.read_data          (io_read_data)                                                                      //                   .export
	);

	nios_system_rs232_0 rs232_0 (
		.clk        (up_clocks_0_sys_clk_clk),                                              //        clock_reset.clk
		.reset      (rst_controller_reset_out_reset),                                       //  clock_reset_reset.reset
		.address    (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address),    // avalon_rs232_slave.address
		.chipselect (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.byteenable (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable), //                   .byteenable
		.read       (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read),       //                   .read
		.write      (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write),      //                   .write
		.writedata  (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.readdata   (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver2_irq),                                             //          interrupt.irq
		.UART_RXD   (rs232_RXD),                                                            // external_interface.export
		.UART_TXD   (rs232_TXD)                                                             //                   .export
	);

	nios_system_pio_0 pio_0 (
		.clk      (up_clocks_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (pio_0_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_0_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (switches_export)                                   // external_connection.export
	);

	nios_system_pio_1 pio_1 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (pio_1_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_1_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_1_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_1_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_1_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (red_leds_export)                                     // external_connection.export
	);

	nios_system_pio_2 pio_2 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                    //               reset.reset_n
		.address    (pio_2_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_2_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_2_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_2_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_2_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (green_leds_export)                                   // external_connection.export
	);

	nios_system_character_lcd_0 character_lcd_0 (
		.clk         (up_clocks_0_sys_clk_clk),                                                     //        clock_reset.clk
		.reset       (rst_controller_reset_out_reset),                                              //  clock_reset_reset.reset
		.address     (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),     //   avalon_lcd_slave.address
		.chipselect  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),  //                   .chipselect
		.read        (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),        //                   .read
		.write       (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),       //                   .write
		.writedata   (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),   //                   .writedata
		.readdata    (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),    //                   .readdata
		.waitrequest (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest), //                   .waitrequest
		.LCD_DATA    (lcd_display_DATA),                                                            // external_interface.export
		.LCD_ON      (lcd_display_ON),                                                              //                   .export
		.LCD_BLON    (lcd_display_BLON),                                                            //                   .export
		.LCD_EN      (lcd_display_EN),                                                              //                   .export
		.LCD_RS      (lcd_display_RS),                                                              //                   .export
		.LCD_RW      (lcd_display_RW)                                                               //                   .export
	);

	nios_system_pio_3 pio_3 (
		.clk      (up_clocks_0_sys_clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (pio_3_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_3_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (push_buttons123_export)                            // external_connection.export
	);

	nios_system_timer_0 timer_0 (
		.clk        (up_clocks_0_sys_clk_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                              //   irq.irq
	);

	nios_system_timer_0 timer_1 (
		.clk        (up_clocks_0_sys_clk_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_1_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_1_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_1_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_1_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_1_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                              //   irq.irq
	);

	nios_system_pio_2 pio_4 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                //               reset.reset_n
		.address    (pio_4_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_4_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_4_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_4_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_4_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex0_1_export)                                       // external_connection.export
	);

	nios_system_pio_2 pio_5 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                //               reset.reset_n
		.address    (pio_5_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_5_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_5_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_5_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_5_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex2_3_export)                                       // external_connection.export
	);

	nios_system_pio_2 pio_6 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                //               reset.reset_n
		.address    (pio_6_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_6_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_6_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_6_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_6_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex4_5_export)                                       // external_connection.export
	);

	nios_system_pio_2 pio_7 (
		.clk        (up_clocks_0_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                //               reset.reset_n
		.address    (pio_7_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_7_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_7_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_7_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_7_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hex6_7_export)                                       // external_connection.export
	);

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),     //                    .address
		.i_avalon_read        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),        //                    .read
		.i_avalon_write       (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),       //                    .write
		.i_avalon_byteenable  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),  //                    .byteenable
		.i_avalon_writedata   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),   //                    .writedata
		.o_avalon_readdata    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),    //                    .readdata
		.o_avalon_waitrequest (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest), //                    .waitrequest
		.i_clock              (up_clocks_0_sys_clk_clk),                                                                             //          clock_sink.clk
		.i_reset_n            (~rst_controller_002_reset_out_reset),                                                                 //    clock_sink_reset.reset_n
		.b_SD_cmd             (sdcard_b_SD_cmd),                                                                                     //         conduit_end.export
		.b_SD_dat             (sdcard_b_SD_dat),                                                                                     //                    .export
		.b_SD_dat3            (sdcard_b_SD_dat3),                                                                                    //                    .export
		.o_SD_clock           (sdcard_o_SD_clock)                                                                                    //                    .export
	);

	amd amd_0 (
		.clk            (up_clocks_0_sys_clk_clk),                                       //          clock.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                           //          reset.reset_n
		.slv_addr       (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_address),   // avalon_slave_0.address
		.slv_start      (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_write),     //               .write
		.slv_data       (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata), //               .writedata
		.slv_done       (),                                                              //               .readyfordata
		.master_wrdata  (amd_0_avalon_master_writedata),                                 //  avalon_master.writedata
		.master_addr    (amd_0_avalon_master_address),                                   //               .address
		.master_rdata   (amd_0_avalon_master_readdata),                                  //               .readdata
		.master_read    (amd_0_avalon_master_read),                                      //               .read
		.master_write   (amd_0_avalon_master_write),                                     //               .write
		.master_waitreq (amd_0_avalon_master_waitrequest)                                //               .waitrequest
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_instruction_master_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                            //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                     //                     reset.reset
		.uav_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (nios2_qsys_0_instruction_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_0_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                               //               (terminated)
		.av_byteenable            (4'b1111),                                                                            //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                                               //               (terminated)
		.av_write                 (1'b0),                                                                               //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                               //               (terminated)
		.av_lock                  (1'b0),                                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                                               //               (terminated)
		.uav_clken                (),                                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                                               //               (terminated)
		.uav_response             (2'b00),                                                                              //               (terminated)
		.av_response              (),                                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_0_data_master_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                     //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                              //                     reset.reset
		.uav_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (nios2_qsys_0_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (nios2_qsys_0_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (nios2_qsys_0_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (nios2_qsys_0_data_master_read),                                               //                          .read
		.av_readdata              (nios2_qsys_0_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (nios2_qsys_0_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (nios2_qsys_0_data_master_write),                                              //                          .write
		.av_writedata             (nios2_qsys_0_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (nios2_qsys_0_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (16),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (2),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (2),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (2),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) amd_0_avalon_master_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                //                       clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                     //                     reset.reset
		.uav_address              (amd_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (amd_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (amd_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (amd_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (amd_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (amd_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (amd_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (amd_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (amd_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (amd_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (amd_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (amd_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (amd_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (amd_0_avalon_master_read),                                               //                          .read
		.av_readdata              (amd_0_avalon_master_readdata),                                           //                          .readdata
		.av_write                 (amd_0_avalon_master_write),                                              //                          .write
		.av_writedata             (amd_0_avalon_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                   //               (terminated)
		.av_byteenable            (2'b11),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                   //               (terminated)
		.av_begintransfer         (1'b0),                                                                   //               (terminated)
		.av_chipselect            (1'b0),                                                                   //               (terminated)
		.av_readdatavalid         (),                                                                       //               (terminated)
		.av_lock                  (1'b0),                                                                   //               (terminated)
		.av_debugaccess           (1'b0),                                                                   //               (terminated)
		.uav_clken                (),                                                                       //               (terminated)
		.av_clken                 (1'b1),                                                                   //               (terminated)
		.uav_response             (2'b00),                                                                  //               (terminated)
		.av_response              (),                                                                       //               (terminated)
		.uav_writeresponserequest (),                                                                       //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                   //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                   //               (terminated)
		.av_writeresponsevalid    ()                                                                        //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_0_jtag_debug_module_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (nios2_qsys_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) new_sdram_controller_0_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                       //                    reset.reset
		.uav_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (new_sdram_controller_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory2_0_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                        //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (onchip_memory2_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (onchip_memory2_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (onchip_memory2_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (onchip_memory2_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken                 (onchip_memory2_0_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read                  (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) to_external_bus_bridge_0_avalon_slave_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                                          //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                                   //                    reset.reset
		.uav_address              (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (to_external_bus_bridge_0_avalon_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                                 //              (terminated)
		.av_lock                  (),                                                                                                 //              (terminated)
		.av_clken                 (),                                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                                 //              (terminated)
		.uav_response             (),                                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) rs232_0_avalon_rs232_slave_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect            (rs232_0_avalon_rs232_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_0_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (pio_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                    //              (terminated)
		.av_read                  (),                                                                    //              (terminated)
		.av_writedata             (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (8),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (1),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (1),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (1),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) character_lcd_0_avalon_lcd_slave_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                                     //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                              //                    reset.reset
		.uav_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (character_lcd_0_avalon_lcd_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                                            //              (terminated)
		.av_burstcount            (),                                                                                            //              (terminated)
		.av_byteenable            (),                                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                                            //              (terminated)
		.av_lock                  (),                                                                                            //              (terminated)
		.av_clken                 (),                                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                                        //              (terminated)
		.av_debugaccess           (),                                                                                            //              (terminated)
		.av_outputenable          (),                                                                                            //              (terminated)
		.uav_response             (),                                                                                            //              (terminated)
		.av_response              (2'b00),                                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_3_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_3_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (pio_3_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                    //              (terminated)
		.av_read                  (),                                                                    //              (terminated)
		.av_writedata             (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_1_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (timer_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (timer_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (timer_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (timer_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (timer_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_4_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_4_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_4_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_4_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_4_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_4_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_5_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_5_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_5_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_5_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_5_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_5_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_6_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_6_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_6_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_6_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_6_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_6_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_7_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_7_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_7_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_7_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_7_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_7_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (8),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                                                  //                    reset.reset
		.uav_address              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                                                    //              (terminated)
		.av_lock                  (),                                                                                                                    //              (terminated)
		.av_clken                 (),                                                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                                                    //              (terminated)
		.uav_response             (),                                                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) amd_0_avalon_slave_0_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                         //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                              //                    reset.reset
		.uav_address              (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_writedata             (amd_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_read                  (),                                                                                //              (terminated)
		.av_readdata              (16'b1101111010101101),                                                            //              (terminated)
		.av_begintransfer         (),                                                                                //              (terminated)
		.av_beginbursttransfer    (),                                                                                //              (terminated)
		.av_burstcount            (),                                                                                //              (terminated)
		.av_byteenable            (),                                                                                //              (terminated)
		.av_readdatavalid         (1'b0),                                                                            //              (terminated)
		.av_waitrequest           (1'b0),                                                                            //              (terminated)
		.av_writebyteenable       (),                                                                                //              (terminated)
		.av_lock                  (),                                                                                //              (terminated)
		.av_chipselect            (),                                                                                //              (terminated)
		.av_clken                 (),                                                                                //              (terminated)
		.uav_clken                (1'b0),                                                                            //              (terminated)
		.av_debugaccess           (),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                //              (terminated)
		.uav_response             (),                                                                                //              (terminated)
		.av_response              (2'b00),                                                                           //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                            //              (terminated)
		.uav_writeresponsevalid   (),                                                                                //              (terminated)
		.av_writeresponserequest  (),                                                                                //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_0_avalon_jtag_slave_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                                         //              (terminated)
		.av_burstcount            (),                                                                                         //              (terminated)
		.av_byteenable            (),                                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                         //              (terminated)
		.av_lock                  (),                                                                                         //              (terminated)
		.av_clken                 (),                                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                                     //              (terminated)
		.av_debugaccess           (),                                                                                         //              (terminated)
		.av_outputenable          (),                                                                                         //              (terminated)
		.uav_response             (),                                                                                         //              (terminated)
		.av_response              (2'b00),                                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_1_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_1_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_1_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_1_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_1_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_1_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_2_s1_translator (
		.clk                      (up_clocks_0_sys_clk_clk),                                             //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pio_2_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pio_2_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (pio_2_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pio_2_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (pio_2_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                    //              (terminated)
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_byteenable            (),                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                     //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.av_address              (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                                       //          .ready
		.av_response             (),                                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_BEGIN_BURST           (87),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.PKT_BURST_TYPE_H          (84),
		.PKT_BURST_TYPE_L          (83),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (99),
		.PKT_THREAD_ID_L           (99),
		.PKT_CACHE_H               (106),
		.PKT_CACHE_L               (103),
		.PKT_DATA_SIDEBAND_H       (86),
		.PKT_DATA_SIDEBAND_L       (86),
		.PKT_QOS_H                 (88),
		.PKT_QOS_L                 (88),
		.PKT_ADDR_SIDEBAND_H       (85),
		.PKT_ADDR_SIDEBAND_L       (85),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                              //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.av_address              (nios2_qsys_0_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (nios2_qsys_0_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (nios2_qsys_0_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                            //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                             //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                            //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_BEGIN_BURST           (69),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_TRANS_EXCLUSIVE       (55),
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_THREAD_ID_H           (81),
		.PKT_THREAD_ID_L           (81),
		.PKT_CACHE_H               (88),
		.PKT_CACHE_L               (85),
		.PKT_DATA_SIDEBAND_H       (68),
		.PKT_DATA_SIDEBAND_L       (68),
		.PKT_QOS_H                 (70),
		.PKT_QOS_L                 (70),
		.PKT_ADDR_SIDEBAND_H       (67),
		.PKT_ADDR_SIDEBAND_L       (67),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.AV_BURSTCOUNT_W           (2),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) amd_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                         //       clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.av_address              (amd_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (amd_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (amd_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (amd_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (amd_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (amd_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (amd_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (amd_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (amd_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (amd_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (amd_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_mux_002_src_valid),                                                      //        rp.valid
		.rp_data                 (rsp_xbar_mux_002_src_data),                                                       //          .data
		.rp_channel              (rsp_xbar_mux_002_src_channel),                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_mux_002_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_mux_002_src_endofpacket),                                                //          .endofpacket
		.rp_ready                (rsp_xbar_mux_002_src_ready),                                                      //          .ready
		.av_response             (),                                                                                // (terminated)
		.av_writeresponserequest (1'b0),                                                                            // (terminated)
		.av_writeresponsevalid   ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                              //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                              //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                               //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                      //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                        //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                            //                .channel
		.rf_sink_ready           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                 //       clk_reset.reset
		.m0_address              (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                                    //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                                    //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                                     //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                              //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                                  //                .channel
		.rf_sink_ready           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                 // clk_reset.reset
		.in_data           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                  //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_002_src_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_mux_002_src_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_mux_002_src_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_mux_002_src_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_002_src_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_mux_002_src_channel),                                                             //                .channel
		.rf_sink_ready           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                  //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                                    //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                             //       clk_reset.reset
		.m0_address              (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                                            //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                                            //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                                             //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                                          //                .channel
		.rf_sink_ready           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                             // clk_reset.reset
		.in_data           (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                                       // (terminated)
		.csr_readdata      (),                                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                       // (terminated)
		.almost_full_data  (),                                                                                                           // (terminated)
		.almost_empty_data (),                                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                                       // (terminated)
		.out_empty         (),                                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                                       // (terminated)
		.out_error         (),                                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                                       // (terminated)
		.out_channel       ()                                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                                    //                .channel
		.rf_sink_ready           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (7),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (60),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_POSTED          (42),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.PKT_TRANS_LOCK            (45),
		.PKT_SRC_ID_H              (66),
		.PKT_SRC_ID_L              (62),
		.PKT_DEST_ID_H             (71),
		.PKT_DEST_ID_L             (67),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (73),
		.PKT_RESPONSE_STATUS_H     (81),
		.PKT_RESPONSE_STATUS_L     (80),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (82),
		.AVS_BURSTCOUNT_W          (1),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                        //       clk_reset.reset
		.m0_address              (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                                       //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                                       //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                                        //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                                               //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                                                 //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                                     //                .channel
		.rf_sink_ready           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (83),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                        // clk_reset.reset
		.in_data           (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                                  // (terminated)
		.csr_readdata      (),                                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                  // (terminated)
		.almost_full_data  (),                                                                                                      // (terminated)
		.almost_empty_data (),                                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                                  // (terminated)
		.out_empty         (),                                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                                  // (terminated)
		.out_error         (),                                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                                  // (terminated)
		.out_channel       ()                                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_3_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_3_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_007_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_007_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_007_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_007_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_007_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_007_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_3_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_3_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_3_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_008_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_008_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_008_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_008_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_008_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_008_src_channel),                                                    //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_009_src_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_mux_009_src_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_mux_009_src_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_mux_009_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_009_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_mux_009_src_channel),                                                    //                .channel
		.rf_sink_ready           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_4_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_4_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_010_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_010_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_010_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_010_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_010_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_010_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_4_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_4_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_4_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_5_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_5_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_011_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_011_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_011_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_011_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_011_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_011_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_5_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_5_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_5_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_6_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_6_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_012_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_012_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_012_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_012_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_012_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_012_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_6_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_6_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_6_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_7_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_7_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_013_src_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_013_src_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_013_src_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_013_src_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_013_src_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_013_src_channel),                                                  //                .channel
		.rf_sink_ready           (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_7_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_7_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_7_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                                            //       clk_reset.reset
		.m0_address              (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_014_src_ready),                                                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_014_src_valid),                                                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_014_src_data),                                                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_014_src_startofpacket),                                                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_014_src_endofpacket),                                                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_014_src_channel),                                                                                                  //                .channel
		.rf_sink_ready           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                                            // clk_reset.reset
		.in_data           (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                                                          // (terminated)
		.csr_readdata      (),                                                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                                          // (terminated)
		.almost_full_data  (),                                                                                                                              // (terminated)
		.almost_empty_data (),                                                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                                                          // (terminated)
		.out_empty         (),                                                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                                                          // (terminated)
		.out_error         (),                                                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                                                          // (terminated)
		.out_channel       ()                                                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (69),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (75),
		.PKT_SRC_ID_L              (71),
		.PKT_DEST_ID_H             (80),
		.PKT_DEST_ID_L             (76),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (84),
		.PKT_PROTECTION_L          (82),
		.PKT_RESPONSE_STATUS_H     (90),
		.PKT_RESPONSE_STATUS_L     (89),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (91),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                   //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                           //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                           //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                            //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                     //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                         //                .channel
		.rf_sink_ready           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                     //     (terminated)
		.m0_writeresponserequest (),                                                                                          //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                       //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (92),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                   //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src16_ready),                                                                     //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src16_valid),                                                                     //                .valid
		.cp_data                 (cmd_xbar_demux_001_src16_data),                                                                      //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src16_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src16_endofpacket),                                                               //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src16_channel),                                                                   //                .channel
		.rf_sink_ready           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                              // (terminated)
		.csr_read          (1'b0),                                                                                               // (terminated)
		.csr_write         (1'b0),                                                                                               // (terminated)
		.csr_readdata      (),                                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                               // (terminated)
		.almost_full_data  (),                                                                                                   // (terminated)
		.almost_empty_data (),                                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                                               // (terminated)
		.out_empty         (),                                                                                                   // (terminated)
		.in_error          (1'b0),                                                                                               // (terminated)
		.out_error         (),                                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                                               // (terminated)
		.out_channel       ()                                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_1_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src17_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src17_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src17_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src17_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src17_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src17_channel),                                              //                .channel
		.rf_sink_ready           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (87),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (89),
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (79),
		.PKT_BURSTWRAP_L           (77),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (102),
		.PKT_PROTECTION_L          (100),
		.PKT_RESPONSE_STATUS_H     (108),
		.PKT_RESPONSE_STATUS_L     (107),
		.PKT_BURST_SIZE_H          (82),
		.PKT_BURST_SIZE_L          (80),
		.ST_CHANNEL_W              (19),
		.ST_DATA_W                 (109),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pio_2_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (up_clocks_0_sys_clk_clk),                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                //       clk_reset.reset
		.m0_address              (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_2_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src18_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src18_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src18_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src18_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src18_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src18_channel),                                              //                .channel
		.rf_sink_ready           (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_2_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (110),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (up_clocks_0_sys_clk_clk),                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.in_data           (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_2_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_2_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	nios_system_addr_router addr_router (
		.sink_ready         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                                       //          .valid
		.src_data           (addr_router_src_data),                                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_system_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios_system_addr_router_002 addr_router_002 (
		.sink_ready         (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (amd_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                       //          .valid
		.src_data           (addr_router_002_src_data),                                                        //          .data
		.src_channel        (addr_router_002_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                  //          .endofpacket
	);

	nios_system_id_router id_router (
		.sink_ready         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                       //       src.ready
		.src_valid          (id_router_src_valid),                                                                       //          .valid
		.src_data           (id_router_src_data),                                                                        //          .data
		.src_channel        (id_router_src_channel),                                                                     //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                               //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                  //          .endofpacket
	);

	nios_system_id_router_001 id_router_001 (
		.sink_ready         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (new_sdram_controller_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                              //       src.ready
		.src_valid          (id_router_001_src_valid),                                                              //          .valid
		.src_data           (id_router_001_src_data),                                                               //          .data
		.src_channel        (id_router_001_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                         //          .endofpacket
	);

	nios_system_id_router id_router_002 (
		.sink_ready         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory2_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                        //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                        //       src.ready
		.src_valid          (id_router_002_src_valid),                                                        //          .valid
		.src_data           (id_router_002_src_data),                                                         //          .data
		.src_channel        (id_router_002_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                   //          .endofpacket
	);

	nios_system_id_router_001 id_router_003 (
		.sink_ready         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (to_external_bus_bridge_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                                          //       src.ready
		.src_valid          (id_router_003_src_valid),                                                                          //          .valid
		.src_data           (id_router_003_src_data),                                                                           //          .data
		.src_channel        (id_router_003_src_channel),                                                                        //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                                  //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                                     //          .endofpacket
	);

	nios_system_id_router id_router_004 (
		.sink_ready         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (rs232_0_avalon_rs232_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                               //       src.ready
		.src_valid          (id_router_004_src_valid),                                                               //          .valid
		.src_data           (id_router_004_src_data),                                                                //          .data
		.src_channel        (id_router_004_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                          //          .endofpacket
	);

	nios_system_id_router id_router_005 (
		.sink_ready         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                             //       src.ready
		.src_valid          (id_router_005_src_valid),                                             //          .valid
		.src_data           (id_router_005_src_data),                                              //          .data
		.src_channel        (id_router_005_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_006 id_router_006 (
		.sink_ready         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (character_lcd_0_avalon_lcd_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                              // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                     //          .valid
		.src_data           (id_router_006_src_data),                                                                      //          .data
		.src_channel        (id_router_006_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                                //          .endofpacket
	);

	nios_system_id_router id_router_007 (
		.sink_ready         (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_3_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                             //       src.ready
		.src_valid          (id_router_007_src_valid),                                             //          .valid
		.src_data           (id_router_007_src_data),                                              //          .data
		.src_channel        (id_router_007_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_008 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                               //          .valid
		.src_data           (id_router_008_src_data),                                                //          .data
		.src_channel        (id_router_008_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                          //          .endofpacket
	);

	nios_system_id_router id_router_009 (
		.sink_ready         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                               //       src.ready
		.src_valid          (id_router_009_src_valid),                                               //          .valid
		.src_data           (id_router_009_src_data),                                                //          .data
		.src_channel        (id_router_009_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                          //          .endofpacket
	);

	nios_system_id_router id_router_010 (
		.sink_ready         (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_4_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                             //       src.ready
		.src_valid          (id_router_010_src_valid),                                             //          .valid
		.src_data           (id_router_010_src_data),                                              //          .data
		.src_channel        (id_router_010_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_011 (
		.sink_ready         (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_5_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                             //       src.ready
		.src_valid          (id_router_011_src_valid),                                             //          .valid
		.src_data           (id_router_011_src_data),                                              //          .data
		.src_channel        (id_router_011_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_012 (
		.sink_ready         (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_6_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                             //       src.ready
		.src_valid          (id_router_012_src_valid),                                             //          .valid
		.src_data           (id_router_012_src_data),                                              //          .data
		.src_channel        (id_router_012_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_013 (
		.sink_ready         (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_7_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                             //       src.ready
		.src_valid          (id_router_013_src_valid),                                             //          .valid
		.src_data           (id_router_013_src_data),                                              //          .data
		.src_channel        (id_router_013_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router id_router_014 (
		.sink_ready         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (altera_up_sd_card_avalon_interface_0_avalon_sdcard_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                                                  // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                                                             //       src.ready
		.src_valid          (id_router_014_src_valid),                                                                                             //          .valid
		.src_data           (id_router_014_src_data),                                                                                              //          .data
		.src_channel        (id_router_014_src_channel),                                                                                           //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                                                                     //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                                                                        //          .endofpacket
	);

	nios_system_id_router_015 id_router_015 (
		.sink_ready         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (amd_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                         //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                                         //       src.ready
		.src_valid          (id_router_015_src_valid),                                                         //          .valid
		.src_data           (id_router_015_src_data),                                                          //          .data
		.src_channel        (id_router_015_src_channel),                                                       //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                                 //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                                    //          .endofpacket
	);

	nios_system_id_router_016 id_router_016 (
		.sink_ready         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                                  //       src.ready
		.src_valid          (id_router_016_src_valid),                                                                  //          .valid
		.src_data           (id_router_016_src_data),                                                                   //          .data
		.src_channel        (id_router_016_src_channel),                                                                //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                             //          .endofpacket
	);

	nios_system_id_router_016 id_router_017 (
		.sink_ready         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                             //       src.ready
		.src_valid          (id_router_017_src_valid),                                             //          .valid
		.src_data           (id_router_017_src_data),                                              //          .data
		.src_channel        (id_router_017_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                        //          .endofpacket
	);

	nios_system_id_router_016 id_router_018 (
		.sink_ready         (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_2_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (up_clocks_0_sys_clk_clk),                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                      // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                             //       src.ready
		.src_valid          (id_router_018_src_valid),                                             //          .valid
		.src_data           (id_router_018_src_data),                                              //          .data
		.src_channel        (id_router_018_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (up_clocks_0_sys_clk_clk),        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (98),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (9),
		.PIPELINED                 (0),
		.ST_DATA_W                 (109),
		.ST_CHANNEL_W              (19),
		.VALID_WIDTH               (19),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (76),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (up_clocks_0_sys_clk_clk),            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter (
		.clk                   (up_clocks_0_sys_clk_clk),             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_001_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_001_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_001_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_001_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_001_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_001_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_001 (
		.clk                   (up_clocks_0_sys_clk_clk),                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (40),
		.PKT_ADDR_L                (9),
		.PKT_BEGIN_BURST           (60),
		.PKT_BYTE_CNT_H            (49),
		.PKT_BYTE_CNT_L            (47),
		.PKT_BYTEEN_H              (8),
		.PKT_BYTEEN_L              (8),
		.PKT_BURST_SIZE_H          (55),
		.PKT_BURST_SIZE_L          (53),
		.PKT_BURST_TYPE_H          (57),
		.PKT_BURST_TYPE_L          (56),
		.PKT_BURSTWRAP_H           (52),
		.PKT_BURSTWRAP_L           (50),
		.PKT_TRANS_COMPRESSED_READ (41),
		.PKT_TRANS_WRITE           (43),
		.PKT_TRANS_READ            (44),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (82),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (47),
		.OUT_BURSTWRAP_H           (52),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_002 (
		.clk                   (up_clocks_0_sys_clk_clk),                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_006_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_006_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_006_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_006_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_006_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_006_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (69),
		.PKT_BYTE_CNT_H            (58),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (64),
		.PKT_BURST_SIZE_L          (62),
		.PKT_BURST_TYPE_H          (66),
		.PKT_BURST_TYPE_L          (65),
		.PKT_BURSTWRAP_H           (61),
		.PKT_BURSTWRAP_L           (59),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (91),
		.ST_CHANNEL_W              (19),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (61),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (3),
		.BURSTWRAP_CONST_VALUE     (3)
	) burst_adapter_003 (
		.clk                   (up_clocks_0_sys_clk_clk),                 //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_015_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_015_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_015_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_015_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_015_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_015_src_ready),              //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (1)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (up_clocks_0_sys_clk_clk),                    //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                             // reset_in0.reset
		.reset_in1  (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk        (clk_clk),                                    //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req  (),                                           // (terminated)
		.reset_in2  (1'b0),                                       // (terminated)
		.reset_in3  (1'b0),                                       // (terminated)
		.reset_in4  (1'b0),                                       // (terminated)
		.reset_in5  (1'b0),                                       // (terminated)
		.reset_in6  (1'b0),                                       // (terminated)
		.reset_in7  (1'b0),                                       // (terminated)
		.reset_in8  (1'b0),                                       // (terminated)
		.reset_in9  (1'b0),                                       // (terminated)
		.reset_in10 (1'b0),                                       // (terminated)
		.reset_in11 (1'b0),                                       // (terminated)
		.reset_in12 (1'b0),                                       // (terminated)
		.reset_in13 (1'b0),                                       // (terminated)
		.reset_in14 (1'b0),                                       // (terminated)
		.reset_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (up_clocks_0_sys_clk_clk),            //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                 (up_clocks_0_sys_clk_clk),            //        clk.clk
		.reset               (rst_controller_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_cmd_src_channel),            //           .channel
		.sink_data           (limiter_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_src15_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (up_clocks_0_sys_clk_clk),                //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket),   //           .endofpacket
		.src14_ready         (cmd_xbar_demux_001_src14_ready),         //      src14.ready
		.src14_valid         (cmd_xbar_demux_001_src14_valid),         //           .valid
		.src14_data          (cmd_xbar_demux_001_src14_data),          //           .data
		.src14_channel       (cmd_xbar_demux_001_src14_channel),       //           .channel
		.src14_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //           .startofpacket
		.src14_endofpacket   (cmd_xbar_demux_001_src14_endofpacket),   //           .endofpacket
		.src15_ready         (cmd_xbar_demux_001_src15_ready),         //      src15.ready
		.src15_valid         (cmd_xbar_demux_001_src15_valid),         //           .valid
		.src15_data          (cmd_xbar_demux_001_src15_data),          //           .data
		.src15_channel       (cmd_xbar_demux_001_src15_channel),       //           .channel
		.src15_startofpacket (cmd_xbar_demux_001_src15_startofpacket), //           .startofpacket
		.src15_endofpacket   (cmd_xbar_demux_001_src15_endofpacket),   //           .endofpacket
		.src16_ready         (cmd_xbar_demux_001_src16_ready),         //      src16.ready
		.src16_valid         (cmd_xbar_demux_001_src16_valid),         //           .valid
		.src16_data          (cmd_xbar_demux_001_src16_data),          //           .data
		.src16_channel       (cmd_xbar_demux_001_src16_channel),       //           .channel
		.src16_startofpacket (cmd_xbar_demux_001_src16_startofpacket), //           .startofpacket
		.src16_endofpacket   (cmd_xbar_demux_001_src16_endofpacket),   //           .endofpacket
		.src17_ready         (cmd_xbar_demux_001_src17_ready),         //      src17.ready
		.src17_valid         (cmd_xbar_demux_001_src17_valid),         //           .valid
		.src17_data          (cmd_xbar_demux_001_src17_data),          //           .data
		.src17_channel       (cmd_xbar_demux_001_src17_channel),       //           .channel
		.src17_startofpacket (cmd_xbar_demux_001_src17_startofpacket), //           .startofpacket
		.src17_endofpacket   (cmd_xbar_demux_001_src17_endofpacket),   //           .endofpacket
		.src18_ready         (cmd_xbar_demux_001_src18_ready),         //      src18.ready
		.src18_valid         (cmd_xbar_demux_001_src18_valid),         //           .valid
		.src18_data          (cmd_xbar_demux_001_src18_data),          //           .data
		.src18_channel       (cmd_xbar_demux_001_src18_channel),       //           .channel
		.src18_startofpacket (cmd_xbar_demux_001_src18_startofpacket), //           .startofpacket
		.src18_endofpacket   (cmd_xbar_demux_001_src18_endofpacket)    //           .endofpacket
	);

	nios_system_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_src_ready),               //     sink0.ready
		.sink0_valid         (width_adapter_src_valid),               //          .valid
		.sink0_channel       (width_adapter_src_channel),             //          .channel
		.sink0_data          (width_adapter_src_data),                //          .data
		.sink0_startofpacket (width_adapter_src_startofpacket),       //          .startofpacket
		.sink0_endofpacket   (width_adapter_src_endofpacket),         //          .endofpacket
		.sink1_ready         (width_adapter_004_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_004_src_valid),           //          .valid
		.sink1_channel       (width_adapter_004_src_channel),         //          .channel
		.sink1_data          (width_adapter_004_src_data),            //          .data
		.sink1_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_002 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src2_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src2_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src2_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src2_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src2_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src2_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_001 cmd_xbar_mux_003 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_001_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_001_src_valid),           //          .valid
		.sink0_channel       (width_adapter_001_src_channel),         //          .channel
		.sink0_data          (width_adapter_001_src_data),            //          .data
		.sink0_startofpacket (width_adapter_001_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_001_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_005_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_005_src_valid),           //          .valid
		.sink1_channel       (width_adapter_005_src_channel),         //          .channel
		.sink1_data          (width_adapter_005_src_data),            //          .data
		.sink1_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_004 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src4_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src4_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src4_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src4_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src4_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src4_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src4_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_005 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src5_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src5_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src5_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src5_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src5_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src5_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src5_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src5_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src5_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src5_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src5_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_006 cmd_xbar_mux_006 (
		.clk                 (up_clocks_0_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_reset_out_reset),      // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_002_src_ready),         //     sink0.ready
		.sink0_valid         (width_adapter_002_src_valid),         //          .valid
		.sink0_channel       (width_adapter_002_src_channel),       //          .channel
		.sink0_data          (width_adapter_002_src_data),          //          .data
		.sink0_startofpacket (width_adapter_002_src_startofpacket), //          .startofpacket
		.sink0_endofpacket   (width_adapter_002_src_endofpacket),   //          .endofpacket
		.sink1_ready         (width_adapter_006_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_006_src_valid),         //          .valid
		.sink1_channel       (width_adapter_006_src_channel),       //          .channel
		.sink1_data          (width_adapter_006_src_data),          //          .data
		.sink1_startofpacket (width_adapter_006_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_006_src_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_007 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src7_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src7_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src7_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src7_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src7_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src7_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src7_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src7_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src7_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src7_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_008 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src8_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src8_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src8_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src8_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src8_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src8_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src8_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src8_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src8_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src8_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src8_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src8_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_009 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src9_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src9_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src9_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src9_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src9_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src9_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src9_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src9_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src9_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src9_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src9_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src9_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_010 (
		.clk                 (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src10_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src10_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src10_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src10_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src10_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src10_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src10_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src10_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src10_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src10_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src10_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_011 (
		.clk                 (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_011_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_011_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_011_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_011_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_011_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_011_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src11_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src11_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src11_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src11_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src11_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src11_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src11_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src11_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src11_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src11_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src11_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_012 (
		.clk                 (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_012_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_012_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_012_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_012_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_012_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_012_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src12_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src12_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src12_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src12_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src12_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src12_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src12_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src12_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src12_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src12_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src12_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_013 (
		.clk                 (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_013_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_013_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_013_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_013_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_013_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_013_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src13_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src13_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src13_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src13_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src13_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src13_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src13_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src13_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src13_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src13_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src13_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux cmd_xbar_mux_014 (
		.clk                 (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),     // clk_reset.reset
		.src_ready           (cmd_xbar_mux_014_src_ready),             //       src.ready
		.src_valid           (cmd_xbar_mux_014_src_valid),             //          .valid
		.src_data            (cmd_xbar_mux_014_src_data),              //          .data
		.src_channel         (cmd_xbar_mux_014_src_channel),           //          .channel
		.src_startofpacket   (cmd_xbar_mux_014_src_startofpacket),     //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_014_src_endofpacket),       //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src14_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src14_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src14_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src14_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src14_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src14_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src14_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src14_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src14_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src14_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src14_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src14_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_mux_015 cmd_xbar_mux_015 (
		.clk                 (up_clocks_0_sys_clk_clk),             //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.src_ready           (cmd_xbar_mux_015_src_ready),          //       src.ready
		.src_valid           (cmd_xbar_mux_015_src_valid),          //          .valid
		.src_data            (cmd_xbar_mux_015_src_data),           //          .data
		.src_channel         (cmd_xbar_mux_015_src_channel),        //          .channel
		.src_startofpacket   (cmd_xbar_mux_015_src_startofpacket),  //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_015_src_endofpacket),    //          .endofpacket
		.sink0_ready         (width_adapter_003_src_ready),         //     sink0.ready
		.sink0_valid         (width_adapter_003_src_valid),         //          .valid
		.sink0_channel       (width_adapter_003_src_channel),       //          .channel
		.sink0_data          (width_adapter_003_src_data),          //          .data
		.sink0_startofpacket (width_adapter_003_src_startofpacket), //          .startofpacket
		.sink0_endofpacket   (width_adapter_003_src_endofpacket),   //          .endofpacket
		.sink1_ready         (width_adapter_007_src_ready),         //     sink1.ready
		.sink1_valid         (width_adapter_007_src_valid),         //          .valid
		.sink1_channel       (width_adapter_007_src_channel),       //          .channel
		.sink1_data          (width_adapter_007_src_data),          //          .data
		.sink1_startofpacket (width_adapter_007_src_startofpacket), //          .startofpacket
		.sink1_endofpacket   (width_adapter_007_src_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (up_clocks_0_sys_clk_clk),           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_001 rsp_xbar_demux_003 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_004 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_005 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_006 rsp_xbar_demux_006 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_007 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_008 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_009 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_010 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_011 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_011_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_011_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_012 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_012_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_012_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_013 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_013_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_013_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux rsp_xbar_demux_014 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_014_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_014_src1_endofpacket)    //          .endofpacket
	);

	nios_system_cmd_xbar_demux_002 rsp_xbar_demux_015 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_015_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_015_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_015_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_015_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_015_src1_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_016 rsp_xbar_demux_016 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_016 rsp_xbar_demux_017 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_demux_016 rsp_xbar_demux_018 (
		.clk                (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid            (rsp_xbar_mux_src_valid),                //          .valid
		.src_data             (rsp_xbar_mux_src_data),                 //          .data
		.src_channel          (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket    (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready          (width_adapter_008_src_ready),           //     sink1.ready
		.sink1_valid          (width_adapter_008_src_valid),           //          .valid
		.sink1_channel        (width_adapter_008_src_channel),         //          .channel
		.sink1_data           (width_adapter_008_src_data),            //          .data
		.sink1_startofpacket  (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket    (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (width_adapter_010_src_ready),           //     sink3.ready
		.sink3_valid          (width_adapter_010_src_valid),           //          .valid
		.sink3_channel        (width_adapter_010_src_channel),         //          .channel
		.sink3_data           (width_adapter_010_src_data),            //          .data
		.sink3_startofpacket  (width_adapter_010_src_startofpacket),   //          .startofpacket
		.sink3_endofpacket    (width_adapter_010_src_endofpacket),     //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (width_adapter_012_src_ready),           //     sink6.ready
		.sink6_valid          (width_adapter_012_src_valid),           //          .valid
		.sink6_channel        (width_adapter_012_src_channel),         //          .channel
		.sink6_data           (width_adapter_012_src_data),            //          .data
		.sink6_startofpacket  (width_adapter_012_src_startofpacket),   //          .startofpacket
		.sink6_endofpacket    (width_adapter_012_src_endofpacket),     //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src0_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink15_ready         (width_adapter_014_src_ready),           //    sink15.ready
		.sink15_valid         (width_adapter_014_src_valid),           //          .valid
		.sink15_channel       (width_adapter_014_src_channel),         //          .channel
		.sink15_data          (width_adapter_014_src_data),            //          .data
		.sink15_startofpacket (width_adapter_014_src_startofpacket),   //          .startofpacket
		.sink15_endofpacket   (width_adapter_014_src_endofpacket)      //          .endofpacket
	);

	nios_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (width_adapter_009_src_ready),           //     sink1.ready
		.sink1_valid          (width_adapter_009_src_valid),           //          .valid
		.sink1_channel        (width_adapter_009_src_channel),         //          .channel
		.sink1_data           (width_adapter_009_src_data),            //          .data
		.sink1_startofpacket  (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket    (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src1_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src1_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink3_ready          (width_adapter_011_src_ready),           //     sink3.ready
		.sink3_valid          (width_adapter_011_src_valid),           //          .valid
		.sink3_channel        (width_adapter_011_src_channel),         //          .channel
		.sink3_data           (width_adapter_011_src_data),            //          .data
		.sink3_startofpacket  (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink3_endofpacket    (width_adapter_011_src_endofpacket),     //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src1_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src1_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src1_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src1_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink6_ready          (width_adapter_013_src_ready),           //     sink6.ready
		.sink6_valid          (width_adapter_013_src_valid),           //          .valid
		.sink6_channel        (width_adapter_013_src_channel),         //          .channel
		.sink6_data           (width_adapter_013_src_data),            //          .data
		.sink6_startofpacket  (width_adapter_013_src_startofpacket),   //          .startofpacket
		.sink6_endofpacket    (width_adapter_013_src_endofpacket),     //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src1_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src1_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src1_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src1_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src1_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src1_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src1_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src1_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src1_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src1_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src1_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src1_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src1_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src1_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src1_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src1_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src1_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src1_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src1_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src1_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src1_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src1_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src1_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src1_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src1_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src1_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src1_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src1_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src1_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src1_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src1_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src1_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src1_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src1_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src1_endofpacket),   //          .endofpacket
		.sink14_ready         (rsp_xbar_demux_014_src1_ready),         //    sink14.ready
		.sink14_valid         (rsp_xbar_demux_014_src1_valid),         //          .valid
		.sink14_channel       (rsp_xbar_demux_014_src1_channel),       //          .channel
		.sink14_data          (rsp_xbar_demux_014_src1_data),          //          .data
		.sink14_startofpacket (rsp_xbar_demux_014_src1_startofpacket), //          .startofpacket
		.sink14_endofpacket   (rsp_xbar_demux_014_src1_endofpacket),   //          .endofpacket
		.sink15_ready         (width_adapter_015_src_ready),           //    sink15.ready
		.sink15_valid         (width_adapter_015_src_valid),           //          .valid
		.sink15_channel       (width_adapter_015_src_channel),         //          .channel
		.sink15_data          (width_adapter_015_src_data),            //          .data
		.sink15_startofpacket (width_adapter_015_src_startofpacket),   //          .startofpacket
		.sink15_endofpacket   (width_adapter_015_src_endofpacket),     //          .endofpacket
		.sink16_ready         (rsp_xbar_demux_016_src0_ready),         //    sink16.ready
		.sink16_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink16_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink16_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.sink16_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink16_endofpacket   (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink17_ready         (rsp_xbar_demux_017_src0_ready),         //    sink17.ready
		.sink17_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink17_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink17_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink17_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink17_endofpacket   (rsp_xbar_demux_017_src0_endofpacket),   //          .endofpacket
		.sink18_ready         (rsp_xbar_demux_018_src0_ready),         //    sink18.ready
		.sink18_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink18_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink18_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink18_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink18_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_system_rsp_xbar_mux_002 rsp_xbar_mux_002 (
		.clk                 (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset               (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src2_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (up_clocks_0_sys_clk_clk),           //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src1_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_001 (
		.clk                  (up_clocks_0_sys_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src3_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src3_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src3_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src3_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src3_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src3_data),            //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (up_clocks_0_sys_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src6_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src6_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src6_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src6_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src6_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src6_data),            //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_003 (
		.clk                  (up_clocks_0_sys_clk_clk),             //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src15_valid),          //      sink.valid
		.in_channel           (cmd_xbar_demux_src15_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_demux_src15_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src15_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_demux_src15_ready),          //          .ready
		.in_data              (cmd_xbar_demux_src15_data),           //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_005 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src3_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src3_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src3_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src3_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (40),
		.OUT_PKT_ADDR_L                (9),
		.OUT_PKT_DATA_H                (7),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (8),
		.OUT_PKT_BYTEEN_L              (8),
		.OUT_PKT_BYTE_CNT_H            (49),
		.OUT_PKT_BYTE_CNT_L            (47),
		.OUT_PKT_TRANS_COMPRESSED_READ (41),
		.OUT_PKT_BURST_SIZE_H          (55),
		.OUT_PKT_BURST_SIZE_L          (53),
		.OUT_PKT_RESPONSE_STATUS_H     (81),
		.OUT_PKT_RESPONSE_STATUS_L     (80),
		.OUT_PKT_TRANS_EXCLUSIVE       (46),
		.OUT_PKT_BURST_TYPE_H          (57),
		.OUT_PKT_BURST_TYPE_L          (56),
		.OUT_ST_DATA_W                 (82),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_006 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src6_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src6_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src6_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src6_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src6_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src6_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (76),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (79),
		.IN_PKT_BURSTWRAP_L            (77),
		.IN_PKT_BURST_SIZE_H           (82),
		.IN_PKT_BURST_SIZE_L           (80),
		.IN_PKT_RESPONSE_STATUS_H      (108),
		.IN_PKT_RESPONSE_STATUS_L      (107),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (84),
		.IN_PKT_BURST_TYPE_L           (83),
		.IN_ST_DATA_W                  (109),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (58),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_BURST_SIZE_H          (64),
		.OUT_PKT_BURST_SIZE_L          (62),
		.OUT_PKT_RESPONSE_STATUS_H     (90),
		.OUT_PKT_RESPONSE_STATUS_L     (89),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_BURST_TYPE_H          (66),
		.OUT_PKT_BURST_TYPE_L          (65),
		.OUT_ST_DATA_W                 (91),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_007 (
		.clk                  (up_clocks_0_sys_clk_clk),                //       clk.clk
		.reset                (rst_controller_reset_out_reset),         // clk_reset.reset
		.in_valid             (cmd_xbar_demux_001_src15_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_001_src15_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_001_src15_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_001_src15_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_001_src15_ready),         //          .ready
		.in_data              (cmd_xbar_demux_001_src15_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_007_src_data),             //          .data
		.out_channel          (width_adapter_007_src_channel),          //          .channel
		.out_valid            (width_adapter_007_src_valid),            //          .valid
		.out_ready            (width_adapter_007_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                                  // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_001_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_001_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_001_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_001_src1_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_010 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src0_data),          //          .data
		.out_endofpacket      (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_010_src_data),            //          .data
		.out_channel          (width_adapter_010_src_channel),         //          .channel
		.out_valid            (width_adapter_010_src_valid),           //          .valid
		.out_ready            (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_010_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_011 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src1_data),          //          .data
		.out_endofpacket      (width_adapter_011_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_011_src_data),            //          .data
		.out_channel          (width_adapter_011_src_channel),         //          .channel
		.out_valid            (width_adapter_011_src_valid),           //          .valid
		.out_ready            (width_adapter_011_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_011_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_012 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_006_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_006_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_006_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_006_src0_data),          //          .data
		.out_endofpacket      (width_adapter_012_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_012_src_data),            //          .data
		.out_channel          (width_adapter_012_src_channel),         //          .channel
		.out_valid            (width_adapter_012_src_valid),           //          .valid
		.out_ready            (width_adapter_012_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_012_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (40),
		.IN_PKT_ADDR_L                 (9),
		.IN_PKT_DATA_H                 (7),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (8),
		.IN_PKT_BYTEEN_L               (8),
		.IN_PKT_BYTE_CNT_H             (49),
		.IN_PKT_BYTE_CNT_L             (47),
		.IN_PKT_TRANS_COMPRESSED_READ  (41),
		.IN_PKT_BURSTWRAP_H            (52),
		.IN_PKT_BURSTWRAP_L            (50),
		.IN_PKT_BURST_SIZE_H           (55),
		.IN_PKT_BURST_SIZE_L           (53),
		.IN_PKT_RESPONSE_STATUS_H      (81),
		.IN_PKT_RESPONSE_STATUS_L      (80),
		.IN_PKT_TRANS_EXCLUSIVE        (46),
		.IN_PKT_BURST_TYPE_H           (57),
		.IN_PKT_BURST_TYPE_L           (56),
		.IN_ST_DATA_W                  (82),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_013 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.in_valid             (rsp_xbar_demux_006_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_006_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_006_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_006_src1_data),          //          .data
		.out_endofpacket      (width_adapter_013_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_013_src_data),            //          .data
		.out_channel          (width_adapter_013_src_channel),         //          .channel
		.out_valid            (width_adapter_013_src_valid),           //          .valid
		.out_ready            (width_adapter_013_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_013_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_014 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_015_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_015_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_015_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_015_src0_data),          //          .data
		.out_endofpacket      (width_adapter_014_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_014_src_data),            //          .data
		.out_channel          (width_adapter_014_src_channel),         //          .channel
		.out_valid            (width_adapter_014_src_valid),           //          .valid
		.out_ready            (width_adapter_014_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_014_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (49),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (58),
		.IN_PKT_BYTE_CNT_L             (56),
		.IN_PKT_TRANS_COMPRESSED_READ  (50),
		.IN_PKT_BURSTWRAP_H            (61),
		.IN_PKT_BURSTWRAP_L            (59),
		.IN_PKT_BURST_SIZE_H           (64),
		.IN_PKT_BURST_SIZE_L           (62),
		.IN_PKT_RESPONSE_STATUS_H      (90),
		.IN_PKT_RESPONSE_STATUS_L      (89),
		.IN_PKT_TRANS_EXCLUSIVE        (55),
		.IN_PKT_BURST_TYPE_H           (66),
		.IN_PKT_BURST_TYPE_L           (65),
		.IN_ST_DATA_W                  (91),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (76),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (82),
		.OUT_PKT_BURST_SIZE_L          (80),
		.OUT_PKT_RESPONSE_STATUS_H     (108),
		.OUT_PKT_RESPONSE_STATUS_L     (107),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (84),
		.OUT_PKT_BURST_TYPE_L          (83),
		.OUT_ST_DATA_W                 (109),
		.ST_CHANNEL_W                  (19),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_015 (
		.clk                  (up_clocks_0_sys_clk_clk),               //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_015_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_015_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_015_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_015_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_015_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_015_src1_data),          //          .data
		.out_endofpacket      (width_adapter_015_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_015_src_data),            //          .data
		.out_channel          (width_adapter_015_src_channel),         //          .channel
		.out_valid            (width_adapter_015_src_valid),           //          .valid
		.out_ready            (width_adapter_015_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_015_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (up_clocks_0_sys_clk_clk),        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

endmodule
